//Celera:switchideal_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU19
//Celera Confidential Symbol Generator
//1000 Ohm pulldownSwitch
module switchideal_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU19 (CELV,O,enable_switch,CELG,CELSUB);
input CELV;
input enable_switch;
inout O;
input CELG;
input CELSUB;
endmodule

