//Celera:delay0_delayfixed_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU30_delay0
//TYPE: fixed 20ns
module delay0_delayfixed_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU30_delay0 (i, CELV, o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELSUB;
input CELG;
endmodule

