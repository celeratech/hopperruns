// ------------------------ Module Definitions -----------
module VESPAasmTIMERminimum_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU11 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU13 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmPRIORITYD2_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU15 (i0,i1,o0,o1,Tstate,CELG59462,CELV96848,CELSUB40948,Tpriority0_0,Tpriority0_1,TpriorityX_0,TpriorityX_1);
  input  i0;
  input  i1;
  output  o0;
  output  o1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  input  Tpriority0_0;
  input  Tpriority0_1;
  input  TpriorityX_0;
  input  TpriorityX_1;
endmodule

module VESPAasmPRIORITYD2_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU18 (i0,i1,o0,o1,Tstate,CELG59462,CELV96848,CELSUB40948,Tpriority0_0,Tpriority0_1,TpriorityX_0,TpriorityX_1);
  input  i0;
  input  i1;
  output  o0;
  output  o1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  input  Tpriority0_0;
  input  Tpriority0_1;
  input  TpriorityX_0;
  input  TpriorityX_1;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU21 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU22 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU23 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU24 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU25 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU26 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR3_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU27 (i0,i1,i2,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR2_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU28 (i0,i1,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU29 (i0,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSTATE4DF_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU3 (r0,r1,s0,s1,porb,state0,state1,state2,state3,CELG59462,CELV96848,hjconfig_0,hjconfig_1,hjconfig_2,CELSUB40948);
  input  r0;
  input  r1;
  input  s0;
  input  s1;
  input  porb;
  output  state0;
  output  state1;
  output  state2;
  output  state3;
  input  CELG59462;
  input  CELV96848;
  input  hjconfig_0;
  input  hjconfig_1;
  input  hjconfig_2;
  input  CELSUB40948;
endmodule

module VESPAasmSR1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU30 (i0,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU31 (o,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU32 (o,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT2_0_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU33 (o,tstate0,tstate1,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate0;
  input  tstate1;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU34 (o,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmTIMERminimum_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU7 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU9 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module inv_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU1 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module oneshot_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU2 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU8 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU10 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU12 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU14 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU35 (i,tdi_SOFTSTARTinternalNOFAULT_OFF,ten_SOFTSTARTinternalNOFAULT_OFF,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_SOFTSTARTinternalNOFAULT_OFF;
  input  ten_SOFTSTARTinternalNOFAULT_OFF;
endmodule

module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU36 (i,tdi_SOFTSTARTinternalNOFAULT_STARTUP,ten_SOFTSTARTinternalNOFAULT_STARTUP,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_SOFTSTARTinternalNOFAULT_STARTUP;
  input  ten_SOFTSTARTinternalNOFAULT_STARTUP;
endmodule

module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU37 (i,tdi_SOFTSTARTinternalNOFAULT_DONE,ten_SOFTSTARTinternalNOFAULT_DONE,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_SOFTSTARTinternalNOFAULT_DONE;
  input  ten_SOFTSTARTinternalNOFAULT_DONE;
endmodule

module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU38 (i,tdi_SOFTSTARTinternalNOFAULT_CHARGE,ten_SOFTSTARTinternalNOFAULT_CHARGE,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_SOFTSTARTinternalNOFAULT_CHARGE;
  input  ten_SOFTSTARTinternalNOFAULT_CHARGE;
endmodule

module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU39 (i,tdi_SOFTSTARTinternalNOFAULT_state_done,ten_SOFTSTARTinternalNOFAULT_state_done,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_SOFTSTARTinternalNOFAULT_state_done;
  input  ten_SOFTSTARTinternalNOFAULT_state_done;
endmodule

module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU40 (i,tdi_SOFTSTARTinternalNOFAULT_state_off,ten_SOFTSTARTinternalNOFAULT_state_off,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_SOFTSTARTinternalNOFAULT_state_off;
  input  ten_SOFTSTARTinternalNOFAULT_state_off;
endmodule

module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU41 (i,tdi_SOFTSTARTinternalNOFAULT_enable_startup,ten_SOFTSTARTinternalNOFAULT_enable_startup,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_SOFTSTARTinternalNOFAULT_enable_startup;
  input  ten_SOFTSTARTinternalNOFAULT_enable_startup;
endmodule

module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU42 (i,tdi_SOFTSTARTinternalNOFAULT_enable_charge,ten_SOFTSTARTinternalNOFAULT_enable_charge,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_SOFTSTARTinternalNOFAULT_enable_charge;
  input  ten_SOFTSTARTinternalNOFAULT_enable_charge;
endmodule

//Verilog HDL for "Generate", "STONEnoconn" "functional"


module STONEnoconn ( noconn );

  input noconn;
endmodule


//Verilog HDL for "DFT", "DFTtm8d" "functional"


module DFTtm8d ( a, ten, tdo, tmi, G, SUB, V, tdi, tma );

  input V;
  input  [7:0] tma;
  output  [7:0] ten;
  output  [1:0] a;
  inout tdo;
  input  [7:0] tdi;
  input G;
  input SUB;
  inout  [4:0] tmi;
endmodule


//Verilog HDL for "DRM", "drm16" "functional"


module drm16 ( V, G, SUB, tmi, bypload, lastdrm, id, por0, por1, drm0, drm1,
d1, d0 );

  input lastdrm;
  input V;
  output d1;
  input  [7:0] id;
  output d0;
  input  [7:0] por1;
  input bypload;
  output  [7:0] drm0;
  input  [7:0] por0;
  input G;
  output  [7:0] drm1;
  inout  [4:0] tmi;
  input SUB;
endmodule


// ------------------------ Module Verilog ---------------
module SOFTSTARTinternalNOFAULT_DYES_XU1_XSTEPDOWN_XSOFTSTART_XU1 (tdo, tmi, porb, CELG59462, CELV96848, state_off, state_done, CELSUB40948, done_measure, enable_charge, ready_startup, enable_startup, enable_softstart);
inout  tdo;
inout [4:0] tmi;
input  porb;
input  CELG59462;
input  CELV96848;
output  state_off;
output  state_done;
input  CELSUB40948;
input  done_measure;
output  enable_charge;
input  ready_startup;
output  enable_startup;
input  enable_softstart;


// ------------------------ Wires ------------------------
wire [4:0] tmi;
wire [1:0] a;
wire [7:0] tdi;
wire [7:0] ten;
wire [7:0] tma;
wire [7:0] id;
wire [7:0] drm0;
wire [7:0] drm1;
wire [7:0] por0;
wire [7:0] por1;

// ------------------------ Networks ---------------------
VESPAasmTIMERminimum_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU11 XU11 (
.state(net_177),
.Tstate(net_190),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_188),
.tmin_delayoutput(net_189)
);

VESPAasmTIMERminimum_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU13 XU13 (
.state(net_164),
.Tstate(net_196),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_192),
.tmin_delayoutput(net_193)
);

VESPAasmPRIORITYD2_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU15 XU15 (
.i0(net_178),
.i1(net_183),
.o0(net_179),
.o1(net_162),
.Tstate(net_174),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.Tpriority0_0(net_117),
.Tpriority0_1(net_118),
.TpriorityX_0(net_119),
.TpriorityX_1(net_120)
);

VESPAasmPRIORITYD2_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU18 XU18 (
.i0(net_194),
.i1(net_195),
.o0(net_168),
.o1(net_175),
.Tstate(net_190),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.Tpriority0_0(net_133),
.Tpriority0_1(net_134),
.TpriorityX_0(net_135),
.TpriorityX_1(net_136)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU21 XU21 (
.o(net_161),
.i0(net_160),
.Tstate(net_167),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU22 XU22 (
.o(net_178),
.i0(ready_startup),
.Tstate(net_174),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU23 XU23 (
.o(net_183),
.i0(net_171),
.Tstate(net_174),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU24 XU24 (
.o(net_191),
.i0(net_171),
.Tstate(net_196),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU25 XU25 (
.o(net_194),
.i0(done_measure),
.Tstate(net_190),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU26 XU26 (
.o(net_195),
.i0(net_171),
.Tstate(net_190),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR3_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU27 XU27 (
.i0(net_162),
.i1(net_168),
.i2(net_175),
.sr(net_163),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR2_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU28 XU28 (
.i0(net_191),
.i1(net_175),
.sr(net_182),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU29 XU29 (
.i0(net_161),
.sr(net_165),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSTATE4DF_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU3 XU3 (
.r0(net_163),
.r1(net_182),
.s0(net_165),
.s1(net_176),
.porb(porb),
.state0(net_159),
.state1(net_166),
.state2(net_164),
.state3(net_177),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.hjconfig_0(net_149),
.hjconfig_1(net_150),
.hjconfig_2(net_151),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR1_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU30 XU30 (
.i0(net_179),
.sr(net_176),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU31 XU31 (
.o(state_done),
.tstate(net_164),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU32 XU32 (
.o(state_off),
.tstate(net_159),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT2_0_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU33 XU33 (
.o(enable_startup),
.tstate0(net_166),
.tstate1(net_177),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU34 XU34 (
.o(enable_charge),
.tstate(net_177),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmTIMERminimum_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU7 XU7 (
.state(net_159),
.Tstate(net_167),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_173),
.tmin_delayoutput(net_172)
);

VESPAasmTIMERminimum_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU9 XU9 (
.state(net_166),
.Tstate(net_174),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_186),
.tmin_delayoutput(net_187)
);

inv_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU1 XU1 (
.i(enable_softstart),
.o(net_171),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

oneshot_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU2 XU2 (
.i(enable_softstart),
.o(net_160),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU8 XU8 (
.i(net_173),
.o(net_172),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU10 XU10 (
.i(net_186),
.o(net_187),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU12 XU12 (
.i(net_188),
.o(net_189),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU14 XU14 (
.i(net_192),
.o(net_193),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU35 XU35 (
.i(net_159),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_SOFTSTARTinternalNOFAULT_OFF(tdi_SOFTSTARTinternalNOFAULT_OFF_XU35),
.ten_SOFTSTARTinternalNOFAULT_OFF(ten_SOFTSTARTinternalNOFAULT_OFF_XU35)
);

dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU36 XU36 (
.i(net_166),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_SOFTSTARTinternalNOFAULT_STARTUP(tdi_SOFTSTARTinternalNOFAULT_STARTUP_XU36),
.ten_SOFTSTARTinternalNOFAULT_STARTUP(ten_SOFTSTARTinternalNOFAULT_STARTUP_XU36)
);

dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU37 XU37 (
.i(net_164),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_SOFTSTARTinternalNOFAULT_DONE(tdi_SOFTSTARTinternalNOFAULT_DONE_XU37),
.ten_SOFTSTARTinternalNOFAULT_DONE(ten_SOFTSTARTinternalNOFAULT_DONE_XU37)
);

dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU38 XU38 (
.i(net_177),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_SOFTSTARTinternalNOFAULT_CHARGE(tdi_SOFTSTARTinternalNOFAULT_CHARGE_XU38),
.ten_SOFTSTARTinternalNOFAULT_CHARGE(ten_SOFTSTARTinternalNOFAULT_CHARGE_XU38)
);

dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU39 XU39 (
.i(state_done),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_SOFTSTARTinternalNOFAULT_state_done(tdi_SOFTSTARTinternalNOFAULT_state_done_XU39),
.ten_SOFTSTARTinternalNOFAULT_state_done(ten_SOFTSTARTinternalNOFAULT_state_done_XU39)
);

dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU40 XU40 (
.i(state_off),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_SOFTSTARTinternalNOFAULT_state_off(tdi_SOFTSTARTinternalNOFAULT_state_off_XU40),
.ten_SOFTSTARTinternalNOFAULT_state_off(ten_SOFTSTARTinternalNOFAULT_state_off_XU40)
);

dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU41 XU41 (
.i(enable_startup),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_SOFTSTARTinternalNOFAULT_enable_startup(tdi_SOFTSTARTinternalNOFAULT_enable_startup_XU41),
.ten_SOFTSTARTinternalNOFAULT_enable_startup(ten_SOFTSTARTinternalNOFAULT_enable_startup_XU41)
);

dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU42 XU42 (
.i(enable_charge),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_SOFTSTARTinternalNOFAULT_enable_charge(tdi_SOFTSTARTinternalNOFAULT_enable_charge_XU42),
.ten_SOFTSTARTinternalNOFAULT_enable_charge(ten_SOFTSTARTinternalNOFAULT_enable_charge_XU42)
);

STONEnoconn XNC152 (
.noconn(net_152)
);

DFTtm8d dft_hex0x23 (
.G(CELG59462),
.V(CELV96848),
.a({a1,a0}),
.SUB(CELSUB40948),
.tdi({tdi_SOFTSTARTinternalNOFAULT_enable_charge_XU42,tdi_SOFTSTARTinternalNOFAULT_enable_startup_XU41,tdi_SOFTSTARTinternalNOFAULT_state_off_XU40,tdi_SOFTSTARTinternalNOFAULT_state_done_XU39,tdi_SOFTSTARTinternalNOFAULT_CHARGE_XU38,tdi_SOFTSTARTinternalNOFAULT_DONE_XU37,tdi_SOFTSTARTinternalNOFAULT_STARTUP_XU36,tdi_SOFTSTARTinternalNOFAULT_OFF_XU35}),
.tdo(tdo),
.ten({ten_SOFTSTARTinternalNOFAULT_enable_charge_XU42,ten_SOFTSTARTinternalNOFAULT_enable_startup_XU41,ten_SOFTSTARTinternalNOFAULT_state_off_XU40,ten_SOFTSTARTinternalNOFAULT_state_done_XU39,ten_SOFTSTARTinternalNOFAULT_CHARGE_XU38,ten_SOFTSTARTinternalNOFAULT_DONE_XU37,ten_SOFTSTARTinternalNOFAULT_STARTUP_XU36,ten_SOFTSTARTinternalNOFAULT_OFF_XU35}),
.tma({a0,a0,a1,a0,a0,a0,a1,a1}),
.tmi(tmi[4:0])
);

drm16 drm_hex0x3a (
.G(CELG59462),
.V(CELV96848),
.d0(c0),
.d1(c1),
.id({c0,c0,c1,c1,c1,c0,c1,c0}),
.SUB(CELSUB40948),
.tmi(tmi[4:0]),
.drm0({net_152,net_151,net_150,net_149,net_136,net_135,net_134,net_133}),
.drm1({noconn_drm16_drm1_7,noconn_drm16_drm1_6,noconn_drm16_drm1_5,noconn_drm16_drm1_4,net_120,net_119,net_118,net_117}),
.por0({c1,c0,c0,c0,c0,c0,c0,c0}),
.por1({c0,c0,c0,c0,c0,c0,c0,c0}),
.bypload(c0),
.lastdrm(c1)
);

STONEnoconn XNCnoconn_drm16_drm1_4 (
.noconn(noconn_drm16_drm1_4)
);

STONEnoconn XNCnoconn_drm16_drm1_5 (
.noconn(noconn_drm16_drm1_5)
);

STONEnoconn XNCnoconn_drm16_drm1_6 (
.noconn(noconn_drm16_drm1_6)
);

STONEnoconn XNCnoconn_drm16_drm1_7 (
.noconn(noconn_drm16_drm1_7)
);

endmodule

