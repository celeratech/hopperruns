//Celera:fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZREP
//Celera Confidential Symbol Generator
//power NMOS:Ron:0.200 Ohm
//Vgs 6V Vds 30V
//Kelvin:yes

module fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZREP (GATE,SOURCE,DRAIN,SOURCEk,DRAINk,IREPLICA,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
inout DRAINk;
inout SOURCEk;
input SUB;
inout IREPLICA;
endmodule

