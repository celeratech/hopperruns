//Celera:inv_XLOOP_XCONTROL_XU33_XU10
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XLOOP_XCONTROL_XU33_XU10 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

