module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU7_XU3 (i,TAI_SOFTSTARToutput,ten_SOFTSTARToutput,CELG,CELSUB,CELV);
input  i;
output  TAI_SOFTSTARToutput;
input  ten_SOFTSTARToutput;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

