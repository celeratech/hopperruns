module dfthijack_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU8 (HJregulationclko,CELG,CELV,CELSUB,ten_HJregulationclkenable,ten_HJregulationclkstatus,HJregulationclk);
output  HJregulationclko;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJregulationclkenable;
input  ten_HJregulationclkstatus;
input  HJregulationclk;
endmodule

