//Celera:switchideal_XLOOP_XDRIVER_XTOPSW_XU11
//Celera Confidential Symbol Generator
//1000 Ohm transmissionSwitch
module switchideal_XLOOP_XDRIVER_XTOPSW_XU11 (CELV,O,I,enable_switchb,CELG,CELSUB);
input CELV;
input I;
input enable_switchb;
inout O;
input CELG;
input CELSUB;
endmodule

