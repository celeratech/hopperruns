//Celera:switchideal_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU8
//Celera Confidential Symbol Generator
//1000 Ohm pullupSwitch
module switchideal_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU8 (CELV,O,enable_switch,CELG,CELSUB);
input CELV;
input enable_switch;
inout O;
input CELG;
input CELSUB;
endmodule

