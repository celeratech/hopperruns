//Celera:fetdriver_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWDRIVER
//Celera Confidential Symbol Generator
//FET DRIVER 'n' Type 0.500 Ron 0.200 Roff 
//Input No Levelshifter
//Gate Sense None
//DFT no
module fetdriver_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWDRIVER (HVPOS,enable_fetdriverhv,global_fetdriver,fetin,GATE,gate_status,
CELG,
SIMPV,
HVNEG,CELSUB); 
input HVPOS;
input enable_fetdriverhv;
input global_fetdriver;
input fetin;
output GATE;
output gate_status;
input SIMPV;
input CELG;
input HVNEG;
input CELSUB;
endmodule

