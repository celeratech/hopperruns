//Celera:switchideal_XLOOP_XREGULATION_XU2_XU17
//Celera Confidential Symbol Generator
//10000 Ohm pulldownSwitch
module switchideal_XLOOP_XREGULATION_XU2_XU17 (CELV,O,enable_switchb,CELG,CELSUB);
input CELV;
input enable_switchb;
inout O;
input CELG;
input CELSUB;
endmodule

