// ------------------------ Module Definitions -----------
// ------------------------ Module Verilog ---------------
module RINGstepdownAugment_XU1_XPADS (EN, SW, OUT, POK, MUDG, MUDV, CBOOT, MUDHV, PMUDG, PMUDV, PMUDHV, sense_OUT, sense_MUDV, kelvin_MUDG);
  input  EN;
  input  SW;
  input  OUT;
  input  POK;
  input  MUDG;
  input  MUDV;
  input  CBOOT;
  input  MUDHV;
  input  PMUDG;
  input  PMUDV;
  input  PMUDHV;
  input  sense_OUT;
  input  sense_MUDV;
  input  kelvin_MUDG;


// ------------------------ Wires ------------------------

// ------------------------ Networks ---------------------
endmodule

