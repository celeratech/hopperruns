//Celera:fet_fet_cboot_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU5_Xnmos_Xfet
//Celera Confidential Symbol Generator
//power NMOS:Ron:10.000 Ohm
//Vgs 6V Vds 40V
//Kelvin:no

module fet_fet_cboot_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU5_Xnmos_Xfet (GATE,SOURCE,DRAIN,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
endmodule

