//Celera:nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU12
//Celera Confidential Symbol Generator
//5V Inverter
module nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU12 (CELV,CELG,i0,i1,i2,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input i2;
input SUB;
output o;
endmodule

