//Celera:inv_XLOOP_XFEEDBACK_XU2_XU18_XU53
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XLOOP_XFEEDBACK_XU2_XU18_XU53 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

