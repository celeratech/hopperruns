//Celera:inv_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU15
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU15 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

