module dftprobe_XLOOP_XREG_XDEBUG_XU6 (i,TAI_REGvc,ten_REGvc,CELG,CELSUB,CELV);
input  i;
output  TAI_REGvc;
input  ten_REGvc;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

