//Celera:amux2_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU20
//Celera Confidential Symbol Generator
//Inputs: 2, Switch On Resistance: 1K
//Type of Control:pin, T-Switch: no
module amux2_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU20 (CELV,SUB,O,I0,I1,
amux,
CELG);
input CELV;
input SUB;
output O;
input I0;
input I1;
input amux;
input CELG;
endmodule

