//Celera:nand4_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU7
//Celera Confidential Symbol Generator
//nand4
module nand4_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU7 (CELV,CELG,i0,i1,i2,i3,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input i2;
input i3;
input SUB;
output o;
endmodule

