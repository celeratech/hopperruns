module dftprobe_XLOOP_XREG_XDEBUG_XU7 (i,tdi_REGgo,ten_REGgo,CELG,CELSUB,CELV);
input  i;
output  tdi_REGgo;
input  ten_REGgo;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

