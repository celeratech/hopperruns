//Celera:dbuf_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU13_XU8
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU13_XU8 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

