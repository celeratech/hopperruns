module dftprobe_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU16 (i,tdi_botswstatus,ten_botswstatus,CELG,CELSUB,CELV);
input  i;
output  tdi_botswstatus;
input  ten_botswstatus;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

