//Celera:dbuf_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU23_XU6
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU23_XU6 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

