module dftprobe_XU1_XSERVICE_XATESERVICE_XU13 (i,tdi_stosc,ten_stosc,CELG,CELSUB,CELV);
input  i;
output  tdi_stosc;
input  ten_stosc;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

