//Celera:inv_XLOOP_XCONTROL_XU64_XU6
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XLOOP_XCONTROL_XU64_XU6 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

