//Celera:tie_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU9
//Celera Confidential Symbol Generator
//TIE
module tie_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU9 (CELV,CELG,a1,SUB);
input CELV;
input CELG;
output a1;
input SUB;
endmodule

