//Celera:nand2_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU12_XU4
//Celera Confidential Symbol Generator
//5V NAND2
module nand2_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU12_XU4 (CELV,CELG,i0,i1,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input SUB;
output o;
endmodule

