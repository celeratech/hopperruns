module dftprobe_XU1_XSERVICE_XATESERVICE_XU8 (i,tdi_stref,ten_stref,CELG,CELSUB,CELV);
input  i;
output  tdi_stref;
input  ten_stref;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

