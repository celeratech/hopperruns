module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU74 (i,tdi_STEPDOWNalgorithmCONTROL0p2_UNDEF5,ten_STEPDOWNalgorithmCONTROL0p2_UNDEF5,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_UNDEF5;
input  ten_STEPDOWNalgorithmCONTROL0p2_UNDEF5;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

