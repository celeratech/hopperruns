//Celera:resistor_resistor_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xpassive
//Celera Confidential Symbol Generator
//RESISTOR:1000.00KOhm TYPE:poly DFT:no
module resistor_resistor_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xpassive (RP,
CELG,
RN);
inout RP;
inout RN;
input CELG;
endmodule

