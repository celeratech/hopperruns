//Celera:decoder3_XLOOP_XCONTROL_XU12_XU13
//Celera Confidential Symbol Generator
//DECODER
module decoder3_XLOOP_XCONTROL_XU12_XU13 (CELV,i,o,
CELG,SUB);
input CELV;
input [2:0] i;
output [7:0] o;
input CELG;
input SUB;
endmodule

