//Celera:dbuf_XLOOP_XDRIVER_XATEDRIVER_XU21
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XLOOP_XDRIVER_XATEDRIVER_XU21 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

