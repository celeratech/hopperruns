module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU79 (i,tdi_STEPDOWNalgorithmCONTROL0p2_fault_control,ten_STEPDOWNalgorithmCONTROL0p2_fault_control,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_fault_control;
input  ten_STEPDOWNalgorithmCONTROL0p2_fault_control;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

