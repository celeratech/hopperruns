module dftprobe_XLOOP_XCONTROL_XU70 (i,tdi_STEPDOWNalgorithmCONTROL1p3_TOP,ten_STEPDOWNalgorithmCONTROL1p3_TOP,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_TOP;
input  ten_STEPDOWNalgorithmCONTROL1p3_TOP;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

