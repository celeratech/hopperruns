//Celera:timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU16
//Celera Confidential Symbol Generator
//TYPE:rise Bits:5 with 2.0ns LSB
module timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU16 (CELV,in,out,
factory_timingskew,
CELG,CELSUB);
input CELV;
input in;
output out;
input [4:0] factory_timingskew;
input CELG;
input CELSUB;
endmodule

