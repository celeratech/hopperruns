module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU12 (i,tdi_STEPDOWNalgorithmCONTROL0p2_top7SYNC,ten_STEPDOWNalgorithmCONTROL0p2_top7SYNC,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_top7SYNC;
input  ten_STEPDOWNalgorithmCONTROL0p2_top7SYNC;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

