//Celera:inv_XLOOP_XDRIVER_XTOPDRIVER_XU33
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XLOOP_XDRIVER_XTOPDRIVER_XU33 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

