//Celera:delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU27
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:fall
module delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU27 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

