//Celera:inv_XU1_XSERVICE_XATESERVICE_XU1_XU15
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSERVICE_XATESERVICE_XU1_XU15 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

