//Celera:thermal
//Celera Confidential Symbol Generator
//Thermal Protector:Rise 140C Fall 120C
 module thermal_XU1_XSERVICE_XREFSERVICE_XU5 (SIMPV,CELBG,IP,enable_thermal,fault_thermal,ten,
CELG,CELSUB);
input SIMPV;
input CELBG;
input IP;
input enable_thermal;
output fault_thermal;
input ten;
input CELG;
input CELSUB;
endmodule

