//Celera:fet_cboot_XLOOP_XDRIVER_XTOPSW_XU21_Xnmos
//Celera Confidential Symbol Generator
//power NMOS:Ron:10.000 Ohm
//Vgs 6V Vds 40V
//Kelvin:no

module fet_cboot_XLOOP_XDRIVER_XTOPSW_XU21_Xnmos (GATE,SOURCE,DRAIN,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
endmodule

