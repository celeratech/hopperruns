//Celera:capacitorfixed_slopecomp_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU9_Xslc
//Celera Confidential Symbol Generator
//CAPACITOR CONTROL:capacitor
//VALUE: 20.00pF TYPE:mim
module capacitorfixed_slopecomp_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU9_Xslc (CP,
CN);
inout CP;
inout CN;
endmodule

