module dftprobe_XU1_XSTEPDOWN_XFAULT_XU1_XU7 (i,tdi_FAULTstartup,ten_FAULTstartup,CELG,CELSUB,CELV);
input  i;
output  tdi_FAULTstartup;
input  ten_FAULTstartup;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

