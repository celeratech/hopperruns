module dfthijack_XLOOP_XDRIVER_XDEBUG_XU21 (HJdrveno,CELG,CELV,CELSUB,ten_HJdrvenenable,ten_HJdrvenstatus,HJdrven);
output  HJdrveno;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJdrvenenable;
input  ten_HJdrvenstatus;
input  HJdrven;
endmodule

