//Celera:logicshifterL2H_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xroffadjust
//Logic Level shifter with Enable
module logicshifterL2H_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xroffadjust (enable_logicshifter,
HVPOS,HVNEG,SIMPV,
in,
out,
CELG,CELSUB);
input HVPOS;
input HVNEG;
input SIMPV;
input [1:0] in;
output [1:0] out;
input enable_logicshifter;
input CELSUB;
input CELG;
endmodule

