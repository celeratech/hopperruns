//Celera:fet_switchideal_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU17_Xnmos0
//Celera Confidential Symbol Generator
//signal NMOS:Ron:10000 Ohm
//Vgs 6V Vds 6V
//Kelvin:no
module fet_switchideal_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU17_Xnmos0 (GATE,SOURCE,DRAIN,NMOSiso6,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
input NMOSiso6;
endmodule

