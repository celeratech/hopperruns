//Celera:delayfixed_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU13_XU14
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:rise
module delayfixed_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU13_XU14 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

