module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU39 (i,tdi_SOFTSTARTinternalNOFAULT_state_done,ten_SOFTSTARTinternalNOFAULT_state_done,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTinternalNOFAULT_state_done;
input  ten_SOFTSTARTinternalNOFAULT_state_done;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

