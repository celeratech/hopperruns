//Celera:inv_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU29
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU29 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

