module dftprobe_XLOOP_XCONTROL_XU73 (i,tdi_STEPDOWNalgorithmCONTROL1p3_fault_controller,ten_STEPDOWNalgorithmCONTROL1p3_fault_controller,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_fault_controller;
input  ten_STEPDOWNalgorithmCONTROL1p3_fault_controller;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

