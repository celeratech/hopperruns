//Celera:tie_XU1_XSTEPDOWN_XCORESTATE_XU32_XU8
//Celera Confidential Symbol Generator
//TIE
module tie_XU1_XSTEPDOWN_XCORESTATE_XU32_XU8 (CELV,CELG,a0,SUB);
input CELV;
input CELG;
output a0;
input SUB;
endmodule

