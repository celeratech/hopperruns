module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU7_XU1 (i,tdi_SOFTSTARTstartup,ten_SOFTSTARTstartup,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTstartup;
input  ten_SOFTSTARTstartup;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

