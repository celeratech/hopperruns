//Celera:tie_XU1_XSTEPDOWN_XCORESTATE_XU38_XU41
//Celera Confidential Symbol Generator
//TIE
module tie_XU1_XSTEPDOWN_XCORESTATE_XU38_XU41 (CELV,CELG,a0,SUB);
input CELV;
input CELG;
output a0;
input SUB;
endmodule

