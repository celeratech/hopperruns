module dfthijack_XU1_XSTEPDOWN_XLOOP_XATE_XU5 (HJclockdrivero,CELG,CELV,CELSUB,ten_HJclockdriverenable,ten_HJclockdriverstatus,HJclockdriver);
output  HJclockdrivero;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJclockdriverenable;
input  ten_HJclockdriverstatus;
input  HJclockdriver;
endmodule

