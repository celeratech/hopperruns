module dfthijack_XLOOP_XFEEDBACK_XDEBUG_XU4 (HIJACKfeedbacko,CELG,CELV,CELSUB,ten_HIJACKfeedbackenable,ten_HIJACKfeedbackstatus,HIJACKfeedback);
output  HIJACKfeedbacko;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HIJACKfeedbackenable;
input  ten_HIJACKfeedbackstatus;
input  HIJACKfeedback;
endmodule

