module dftprobe_XLOOP_XDRIVER_XDEBUG_XU15 (i,tdi_DRVbotswipeak,ten_DRVbotswipeak,CELG,CELSUB,CELV);
input  i;
output  tdi_DRVbotswipeak;
input  ten_DRVbotswipeak;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

