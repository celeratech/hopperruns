module dftprobe_XLOOP_XCONTROL_XU68 (i,tdi_STEPDOWNalgorithmCONTROL1p3_UNDEF5,ten_STEPDOWNalgorithmCONTROL1p3_UNDEF5,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_UNDEF5;
input  ten_STEPDOWNalgorithmCONTROL1p3_UNDEF5;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

