module dftprobe_XU1_XSTEPDOWN_XDISCHARGE_XU4_XU2 (i,tdi_DISCHARGEtime,ten_DISCHARGEtime,CELG,CELSUB,CELV);
input  i;
output  tdi_DISCHARGEtime;
input  ten_DISCHARGEtime;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

