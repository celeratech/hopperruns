module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU81 (i,tdi_STEPDOWNalgorithmCORE0p0_UNDEF5,ten_STEPDOWNalgorithmCORE0p0_UNDEF5,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_UNDEF5;
input  ten_STEPDOWNalgorithmCORE0p0_UNDEF5;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

