//Celera:delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU8
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:rise
module delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU8 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

