//Celera:nand2_XLOOP_XDRIVER_XBBM_XU16
//Celera Confidential Symbol Generator
//5V NAND2
module nand2_XLOOP_XDRIVER_XBBM_XU16 (CELV,CELG,i0,i1,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input SUB;
output o;
endmodule

