//Celera:delay0_pulsestretch_XU1_XSTEPDOWN_XFAULT_XU6_XU3_Xpulse
//TYPE: fixed 10ns
module delay0_pulsestretch_XU1_XSTEPDOWN_XFAULT_XU6_XU3_Xpulse (i, CELV, o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELSUB;
input CELG;
endmodule

