module dfthijack_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU6 (hjbotstateo,CELG,CELV,CELSUB,ten_hjbotstateenable,ten_hjbotstatestatus,hjbotstate);
output  hjbotstateo;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_hjbotstateenable;
input  ten_hjbotstatestatus;
input  hjbotstate;
endmodule

