//Celera:fet_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWDRIVER_Xnmos0
//Celera Confidential Symbol Generator
//power NMOS:Ron:1.000 Ohm
//Vgs 6V Vds 6V
//Kelvin:no

module fet_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWDRIVER_Xnmos0 (GATE,SOURCE,DRAIN,NMOSiso6,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
input NMOSiso6;
endmodule

