//Celera:cboot_XLOOP_XDRIVER_XTOPDRIVER_XU5
//Celera Confidential Symbol Generator
//Input: 6V Output: 36CBOOT:Ron:10 Ohm
//Vgs 6V
 //OK Output:low_voltage
module cboot_XLOOP_XDRIVER_XTOPDRIVER_XU5 (CBOOT,SIMPV,CELPOS,on_highside,global_cboot,enable_cboot,ok_cbootlv,SWITCH,CELG,CELSUB);
input CBOOT;
input SWITCH;
input SIMPV;
input CELPOS;
input global_cboot;
input enable_cboot;
input on_highside;
output ok_cbootlv;
input CELG;
input CELSUB;
endmodule

