module dftprobe_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU24 (i,tdi_driverstartup,ten_driverstartup,CELG,CELSUB,CELV);
input  i;
output  tdi_driverstartup;
input  ten_driverstartup;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

