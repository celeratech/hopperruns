module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU73 (i,tdi_STEPDOWNalgorithmCONTROL0p2_UNDEF4,ten_STEPDOWNalgorithmCONTROL0p2_UNDEF4,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_UNDEF4;
input  ten_STEPDOWNalgorithmCONTROL0p2_UNDEF4;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

