//Celera:delay0_delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU31_XU3_delay0
//TYPE: fixed 1ns
module delay0_delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU31_XU3_delay0 (i, CELV, o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELSUB;
input CELG;
endmodule

