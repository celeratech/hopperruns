module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU91 (i,tdi_STEPDOWNalgorithmCORE0p0_fault_core,ten_STEPDOWNalgorithmCORE0p0_fault_core,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_fault_core;
input  ten_STEPDOWNalgorithmCORE0p0_fault_core;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

