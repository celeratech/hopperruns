//Celera:resistor_XLOOP_XREGULATION_XU2_XU34
//Celera Confidential Symbol Generator
//RESISTOR:1000KOhm TYPE:poly DFT:no
module resistor_XLOOP_XREGULATION_XU2_XU34 (RP,
CELG,
RN);
inout RP;
inout RN;
input CELG;
endmodule

