//Celera:resistordivider_vbias_XU1_XSERVICE_XBIASSERVICE_XU1_XRfeedback
//Celera Confidential Symbol Generator
//VMAX:6V R:5000.0KOhm 1Taps
module resistordivider_vbias_XU1_XSERVICE_XBIASSERVICE_XU1_XRfeedback (TOP,
TAP0,
CELG, BOTTOM);
inout TOP;
output TAP0;
input CELG;
inout BOTTOM;
endmodule

