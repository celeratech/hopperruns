module dftprobe_XLOOP_XDRIVER_XDEBUG_XU16 (i,tdi_DRVbotswstatus,ten_DRVbotswstatus,CELG,CELSUB,CELV);
input  i;
output  tdi_DRVbotswstatus;
input  ten_DRVbotswstatus;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

