module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU87 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_softstart,ten_STEPDOWNalgorithmCORE0p0_enable_softstart,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_enable_softstart;
input  ten_STEPDOWNalgorithmCORE0p0_enable_softstart;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

