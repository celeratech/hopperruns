//Celera:delayfixed_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU9_XU30
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:rise
module delayfixed_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU9_XU30 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

