//Celera:dbuf_XLOOP_XDRIVER_XBBM_XU12
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XLOOP_XDRIVER_XBBM_XU12 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

