//Celera:delay0_delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU12_delay0
//TYPE: fixed 100ns
module delay0_delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU12_delay0 (i, CELV, o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELSUB;
input CELG;
endmodule

