//Celera:tie_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU15_XU8
//Celera Confidential Symbol Generator
//TIE
module tie_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU15_XU8 (CELV,CELG,a0,SUB);
input CELV;
input CELG;
output a0;
input SUB;
endmodule

