//Celera:dbuf_XU1_XSTEPDOWN_XFAULT_XU6_XU11
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XFAULT_XU6_XU11 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

