//Celera:switchideal_XLOOP_XREGULATION_XU2_XU11
//Celera Confidential Symbol Generator
//1000 Ohm gndSwitch
module switchideal_XLOOP_XREGULATION_XU2_XU11 (CELV,O,I,enable_switch,CELG,CELSUB);
input CELV;
input I;
input enable_switch;
inout O;
input CELG;
input CELSUB;
endmodule

