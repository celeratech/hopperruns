module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU10 (i,tdi_STEPDOWNalgorithmCONTROL0p2_top1SYNC,ten_STEPDOWNalgorithmCONTROL0p2_top1SYNC,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_top1SYNC;
input  ten_STEPDOWNalgorithmCONTROL0p2_top1SYNC;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

