//Celera:dbuf_XLOOP_XDRIVER_XDEBUG_XU24
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XLOOP_XDRIVER_XDEBUG_XU24 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

