module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU14 (i,tdi_STEPDOWNalgorithmCONTROL0p2_top6SYNC,ten_STEPDOWNalgorithmCONTROL0p2_top6SYNC,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_top6SYNC;
input  ten_STEPDOWNalgorithmCONTROL0p2_top6SYNC;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

