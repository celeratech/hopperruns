//Celera:resistor_resistor_fetdriver_XLOOP_XDRIVER_XBOTSW_XU3_Xpassive
//Celera Confidential Symbol Generator
//RESISTOR:1000.00KOhm TYPE:poly DFT:no
module resistor_resistor_fetdriver_XLOOP_XDRIVER_XBOTSW_XU3_Xpassive (RP,
CELG,
RN);
inout RP;
inout RN;
input CELG;
endmodule

