// ------------------------ Module Definitions -----------
module VESPAclockSYNC_XLOOP_XCONTROL_XU10 (din,out,clock,state,CELG59462,CELV96848,CELSUB40948);
  input  din;
  output  out;
  input  clock;
  input  state;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSTATE8PS_XLOOP_XCONTROL_XU11 (r0,r1,r2,s0,s1,s2,porb,state0,state1,state2,state3,state4,state5,state6,state7,CELG59462,CELV96848,CELSUB40948);
  input  r0;
  input  r1;
  input  r2;
  input  s0;
  input  s1;
  input  s2;
  input  porb;
  output  state0;
  output  state1;
  output  state2;
  output  state3;
  output  state4;
  output  state5;
  output  state6;
  output  state7;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU12 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XLOOP_XCONTROL_XU14 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU17 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU19 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU21 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XLOOP_XCONTROL_XU23 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU26 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XLOOP_XCONTROL_XU28 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmPRIORITY3_XLOOP_XCONTROL_XU31 (i0,i1,i2,o0,o1,o2,Tstate,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  o0;
  output  o1;
  output  o2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmPRIORITY2_XLOOP_XCONTROL_XU32 (i0,i1,o0,o1,Tstate,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  o0;
  output  o1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmPRIORITY2_XLOOP_XCONTROL_XU33 (i0,i1,o0,o1,Tstate,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  o0;
  output  o1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmPRIORITY5_XLOOP_XCONTROL_XU34 (i0,i1,i2,i3,i4,o0,o1,o2,o3,o4,Tstate,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  output  o0;
  output  o1;
  output  o2;
  output  o3;
  output  o4;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmPRIORITY3_XLOOP_XCONTROL_XU35 (i0,i1,i2,o0,o1,o2,Tstate,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  o0;
  output  o1;
  output  o2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU36 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT2_XLOOP_XCONTROL_XU37 (o,i0,i1,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU38 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU39 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU40 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT4_XLOOP_XCONTROL_XU41 (o,i0,i1,i2,i3,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU42 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT4_XLOOP_XCONTROL_XU43 (o,i0,i1,i2,i3,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU44 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU45 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT5_XLOOP_XCONTROL_XU46 (o,i0,i1,i2,i3,i4,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT4_XLOOP_XCONTROL_XU47 (o,i0,i1,i2,i3,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT4_XLOOP_XCONTROL_XU48 (o,i0,i1,i2,i3,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT3_XLOOP_XCONTROL_XU49 (o,i0,i1,i2,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU50 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT2_XLOOP_XCONTROL_XU51 (o,i0,i1,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT2_XLOOP_XCONTROL_XU52 (o,i0,i1,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU53 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR7_XLOOP_XCONTROL_XU54 (i0,i1,i2,i3,i4,i5,i6,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  input  i5;
  input  i6;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR6_XLOOP_XCONTROL_XU55 (i0,i1,i2,i3,i4,i5,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  input  i5;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR3_XLOOP_XCONTROL_XU56 (i0,i1,i2,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR3_XLOOP_XCONTROL_XU57 (i0,i1,i2,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR4_XLOOP_XCONTROL_XU58 (i0,i1,i2,i3,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR1_XLOOP_XCONTROL_XU59 (i0,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_0_XLOOP_XCONTROL_XU60 (o,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT2_0_XLOOP_XCONTROL_XU61 (o,tstate0,tstate1,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate0;
  input  tstate1;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_0_XLOOP_XCONTROL_XU62 (o,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAclocktree3_XLOOP_XCONTROL_XU7 (clock0,clock1,clock2,clocki,CELG59462,CELV96848,CELSUB40948);
  output  clock0;
  output  clock1;
  output  clock2;
  input  clocki;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAclockSYNC_XLOOP_XCONTROL_XU8 (din,out,clock,state,CELG59462,CELV96848,CELSUB40948);
  input  din;
  output  out;
  input  clock;
  input  state;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAclockSYNC_XLOOP_XCONTROL_XU9 (din,out,clock,state,CELG59462,CELV96848,CELSUB40948);
  input  din;
  output  out;
  input  clock;
  input  state;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module inv_XLOOP_XCONTROL_XU1 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU2 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU3 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU4 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU5 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU6 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module delayfixed_XLOOP_XCONTROL_XU13 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU15 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU16 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU18 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU20 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU22 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU24 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU25 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU27 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU29 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU30 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module dftprobe_XLOOP_XCONTROL_XU63 (i,tdi_STEPDOWNalgorithmCONTROL1p3_OFF,ten_STEPDOWNalgorithmCONTROL1p3_OFF,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_OFF;
  input  ten_STEPDOWNalgorithmCONTROL1p3_OFF;
endmodule

module dftprobe_XLOOP_XCONTROL_XU64 (i,tdi_STEPDOWNalgorithmCONTROL1p3_POWERUP,ten_STEPDOWNalgorithmCONTROL1p3_POWERUP,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_POWERUP;
  input  ten_STEPDOWNalgorithmCONTROL1p3_POWERUP;
endmodule

module dftprobe_XLOOP_XCONTROL_XU65 (i,tdi_STEPDOWNalgorithmCONTROL1p3_FAULT,ten_STEPDOWNalgorithmCONTROL1p3_FAULT,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_FAULT;
  input  ten_STEPDOWNalgorithmCONTROL1p3_FAULT;
endmodule

module dftprobe_XLOOP_XCONTROL_XU66 (i,tdi_STEPDOWNalgorithmCONTROL1p3_READY,ten_STEPDOWNalgorithmCONTROL1p3_READY,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_READY;
  input  ten_STEPDOWNalgorithmCONTROL1p3_READY;
endmodule

module dftprobe_XLOOP_XCONTROL_XU67 (i,tdi_STEPDOWNalgorithmCONTROL1p3_IDLE,ten_STEPDOWNalgorithmCONTROL1p3_IDLE,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_IDLE;
  input  ten_STEPDOWNalgorithmCONTROL1p3_IDLE;
endmodule

module dftprobe_XLOOP_XCONTROL_XU68 (i,tdi_STEPDOWNalgorithmCONTROL1p3_UNDEF5,ten_STEPDOWNalgorithmCONTROL1p3_UNDEF5,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_UNDEF5;
  input  ten_STEPDOWNalgorithmCONTROL1p3_UNDEF5;
endmodule

module dftprobe_XLOOP_XCONTROL_XU69 (i,tdi_STEPDOWNalgorithmCONTROL1p3_BOTTOM,ten_STEPDOWNalgorithmCONTROL1p3_BOTTOM,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_BOTTOM;
  input  ten_STEPDOWNalgorithmCONTROL1p3_BOTTOM;
endmodule

module dftprobe_XLOOP_XCONTROL_XU70 (i,tdi_STEPDOWNalgorithmCONTROL1p3_TOP,ten_STEPDOWNalgorithmCONTROL1p3_TOP,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_TOP;
  input  ten_STEPDOWNalgorithmCONTROL1p3_TOP;
endmodule

module dftprobe_XLOOP_XCONTROL_XU71 (i,tdi_STEPDOWNalgorithmCONTROL1p3_topstate,ten_STEPDOWNalgorithmCONTROL1p3_topstate,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_topstate;
  input  ten_STEPDOWNalgorithmCONTROL1p3_topstate;
endmodule

module dftprobe_XLOOP_XCONTROL_XU72 (i,tdi_STEPDOWNalgorithmCONTROL1p3_botstate,ten_STEPDOWNalgorithmCONTROL1p3_botstate,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_botstate;
  input  ten_STEPDOWNalgorithmCONTROL1p3_botstate;
endmodule

module dftprobe_XLOOP_XCONTROL_XU73 (i,tdi_STEPDOWNalgorithmCONTROL1p3_fault_controller,ten_STEPDOWNalgorithmCONTROL1p3_fault_controller,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCONTROL1p3_fault_controller;
  input  ten_STEPDOWNalgorithmCONTROL1p3_fault_controller;
endmodule

//Verilog HDL for "DFT", "DFTtm8d" "functional"


module DFTtm8d ( a, ten, tdo, tmi, G, SUB, V, tdi, tma );

  input V;
  input  [7:0] tma;
  output  [7:0] ten;
  output  [1:0] a;
  inout tdo;
  input  [7:0] tdi;
  input G;
  input SUB;
  inout  [4:0] tmi;
endmodule


//Verilog HDL for "Generate", "STONEnoconn" "functional"


module STONEnoconn ( noconn );

  input noconn;
endmodule


// ------------------------ Module Verilog ---------------
module DRIVERaugment0CONTROL1p_XLOOP_XCONTROL (tdo, tmi, porb, clock, botstate, topstate, CELG59462, CELV96848, go_driver, ok_driver, botswipeak, topswipeak, CELSUB40948, botswzcross, enable_control, freeze_control, switch_control, fault_controller);
inout  tdo;
input [4:0] tmi;
input  porb;
input  clock;
output  botstate;
output  topstate;
input  CELG59462;
input  CELV96848;
input  go_driver;
input  ok_driver;
input  botswipeak;
input  topswipeak;
input  CELSUB40948;
input  botswzcross;
input  enable_control;
input  freeze_control;
input  switch_control;
output  fault_controller;


// ------------------------ Wires ------------------------
wire [4:0] tmi;
wire [1:0] a;
wire [7:0] tdi;
wire [7:0] ten;
wire [7:0] tma;

// ------------------------ Networks ---------------------
VESPAclockSYNC_XLOOP_XCONTROL_XU10 XU10 (
.din(net_346),
.out(net_347),
.clock(net_310),
.state(net_331),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSTATE8PS_XLOOP_XCONTROL_XU11 XU11 (
.r0(net_299),
.r1(net_321),
.r2(net_330),
.s0(net_302),
.s1(net_317),
.s2(net_324),
.porb(porb),
.state0(net_294),
.state1(net_303),
.state2(net_312),
.state3(net_311),
.state4(net_322),
.state5(net_325),
.state6(net_331),
.state7(net_300),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU12 XU12 (
.state(net_294),
.Tstate(net_304),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_314),
.tmin_delayoutput(net_313)
);

VESPAasmTIMERminmax_XLOOP_XCONTROL_XU14 XU14 (
.state(net_303),
.Tstate(net_295),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_338),
.t_delayinput(net_335),
.tmax_delayoutput(net_339),
.tmin_delayoutput(net_336)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU17 XU17 (
.state(net_312),
.Tstate(net_343),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_349),
.tmin_delayoutput(net_348)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU19 XU19 (
.state(net_311),
.Tstate(net_350),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_361),
.tmin_delayoutput(net_360)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU21 XU21 (
.state(net_322),
.Tstate(net_363),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_365),
.tmin_delayoutput(net_364)
);

VESPAasmTIMERminmax_XLOOP_XCONTROL_XU23 XU23 (
.state(net_325),
.Tstate(net_369),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_371),
.t_delayinput(net_372),
.tmax_delayoutput(net_373),
.tmin_delayoutput(net_370)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU26 XU26 (
.state(net_331),
.Tstate(net_374),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_376),
.tmin_delayoutput(net_375)
);

VESPAasmTIMERminmax_XLOOP_XCONTROL_XU28 XU28 (
.state(net_300),
.Tstate(net_377),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_380),
.t_delayinput(net_383),
.tmax_delayoutput(net_382),
.tmin_delayoutput(net_379)
);

VESPAasmPRIORITY3_XLOOP_XCONTROL_XU31 XU31 (
.i0(net_305),
.i1(net_315),
.i2(net_318),
.o0(net_306),
.o1(net_298),
.o2(net_307),
.Tstate(net_295),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmPRIORITY2_XLOOP_XCONTROL_XU32 XU32 (
.i0(net_293),
.i1(net_353),
.o0(net_352),
.o1(net_316),
.Tstate(net_350),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmPRIORITY2_XLOOP_XCONTROL_XU33 XU33 (
.i0(net_334),
.i1(net_368),
.o0(net_367),
.o1(net_366),
.Tstate(net_363),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmPRIORITY5_XLOOP_XCONTROL_XU34 XU34 (
.i0(net_347),
.i1(net_381),
.i2(net_384),
.i3(net_385),
.i4(net_386),
.o0(net_378),
.o1(net_354),
.o2(net_355),
.o3(net_358),
.o4(net_359),
.Tstate(net_374),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmPRIORITY3_XLOOP_XCONTROL_XU35 XU35 (
.i0(net_387),
.i1(net_388),
.i2(net_389),
.o0(net_323),
.o1(net_326),
.o2(net_332),
.Tstate(net_377),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU36 XU36 (
.o(net_297),
.i0(enable_control),
.Tstate(net_304),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT2_XLOOP_XCONTROL_XU37 XU37 (
.o(net_305),
.i0(clock),
.i1(ok_driver),
.Tstate(net_295),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU38 XU38 (
.o(net_315),
.i0(net_338),
.Tstate(net_295),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU39 XU39 (
.o(net_318),
.i0(net_309),
.Tstate(net_295),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU40 XU40 (
.o(net_351),
.i0(net_309),
.Tstate(net_343),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT4_XLOOP_XCONTROL_XU41 XU41 (
.o(net_292),
.i0(go_driver),
.i1(switch_control),
.i2(clock),
.i3(net_329),
.Tstate(net_350),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU42 XU42 (
.o(net_353),
.i0(net_309),
.Tstate(net_350),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT4_XLOOP_XCONTROL_XU43 XU43 (
.o(net_333),
.i0(clock),
.i1(go_driver),
.i2(net_329),
.i3(switch_control),
.Tstate(net_363),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU44 XU44 (
.o(net_368),
.i0(net_309),
.Tstate(net_363),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU45 XU45 (
.o(net_319),
.i0(net_371),
.Tstate(net_369),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT5_XLOOP_XCONTROL_XU46 XU46 (
.o(net_346),
.i0(net_341),
.i1(clock),
.i2(go_driver),
.i3(net_329),
.i4(switch_control),
.Tstate(net_374),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT4_XLOOP_XCONTROL_XU47 XU47 (
.o(net_381),
.i0(botswzcross),
.i1(clock),
.i2(go_driver),
.i3(net_329),
.Tstate(net_374),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT4_XLOOP_XCONTROL_XU48 XU48 (
.o(net_384),
.i0(net_341),
.i1(botswzcross),
.i2(net_345),
.i3(net_329),
.Tstate(net_374),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT3_XLOOP_XCONTROL_XU49 XU49 (
.o(net_385),
.i0(freeze_control),
.i1(clock),
.i2(go_driver),
.Tstate(net_374),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU50 XU50 (
.o(net_386),
.i0(net_309),
.Tstate(net_374),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT2_XLOOP_XCONTROL_XU51 XU51 (
.o(net_387),
.i0(topswipeak),
.i1(clock),
.Tstate(net_377),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT2_XLOOP_XCONTROL_XU52 XU52 (
.o(net_388),
.i0(net_357),
.i1(net_362),
.Tstate(net_377),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU53 XU53 (
.o(net_389),
.i0(net_380),
.Tstate(net_377),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR7_XLOOP_XCONTROL_XU54 XU54 (
.i0(net_298),
.i1(net_307),
.i2(net_316),
.i3(net_319),
.i4(net_323),
.i5(net_326),
.i6(net_332),
.sr(net_299),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR6_XLOOP_XCONTROL_XU55 XU55 (
.i0(net_351),
.i1(net_316),
.i2(net_354),
.i3(net_355),
.i4(net_358),
.i5(net_359),
.sr(net_321),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR3_XLOOP_XCONTROL_XU56 XU56 (
.i0(net_366),
.i1(net_319),
.i2(net_359),
.sr(net_330),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR3_XLOOP_XCONTROL_XU57 XU57 (
.i0(net_297),
.i1(net_367),
.i2(net_378),
.sr(net_302),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR4_XLOOP_XCONTROL_XU58 XU58 (
.i0(net_306),
.i1(net_298),
.i2(net_367),
.i3(net_319),
.sr(net_317),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR1_XLOOP_XCONTROL_XU59 XU59 (
.i0(net_352),
.sr(net_324),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_0_XLOOP_XCONTROL_XU60 XU60 (
.o(topstate),
.tstate(net_300),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT2_0_XLOOP_XCONTROL_XU61 XU61 (
.o(botstate),
.tstate0(net_331),
.tstate1(net_303),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_0_XLOOP_XCONTROL_XU62 XU62 (
.o(fault_controller),
.tstate(net_312),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAclocktree3_XLOOP_XCONTROL_XU7 XU7 (
.clock0(net_291),
.clock1(net_301),
.clock2(net_310),
.clocki(clock),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAclockSYNC_XLOOP_XCONTROL_XU8 XU8 (
.din(net_292),
.out(net_293),
.clock(net_291),
.state(net_311),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAclockSYNC_XLOOP_XCONTROL_XU9 XU9 (
.din(net_333),
.out(net_334),
.clock(net_301),
.state(net_322),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

inv_XLOOP_XCONTROL_XU1 XU1 (
.i(enable_control),
.o(net_309),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU2 XU2 (
.i(freeze_control),
.o(net_329),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU3 XU3 (
.i(botswipeak),
.o(net_341),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU4 XU4 (
.i(go_driver),
.o(net_345),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU5 XU5 (
.i(topswipeak),
.o(net_357),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU6 XU6 (
.i(clock),
.o(net_362),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

delayfixed_XLOOP_XCONTROL_XU13 XU13 (
.i(net_314),
.o(net_313),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU15 XU15 (
.i(net_335),
.o(net_336),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU16 XU16 (
.i(net_335),
.o(net_339),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU18 XU18 (
.i(net_349),
.o(net_348),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU20 XU20 (
.i(net_361),
.o(net_360),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU22 XU22 (
.i(net_365),
.o(net_364),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU24 XU24 (
.i(net_372),
.o(net_370),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU25 XU25 (
.i(net_372),
.o(net_373),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU27 XU27 (
.i(net_376),
.o(net_375),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU29 XU29 (
.i(net_383),
.o(net_379),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU30 XU30 (
.i(net_383),
.o(net_382),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

dftprobe_XLOOP_XCONTROL_XU63 XU63 (
.i(net_294),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_OFF(tdi_STEPDOWNalgorithmCONTROL1p3_OFF_XU63),
.ten_STEPDOWNalgorithmCONTROL1p3_OFF(ten_STEPDOWNalgorithmCONTROL1p3_OFF_XU63)
);

dftprobe_XLOOP_XCONTROL_XU64 XU64 (
.i(net_303),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_POWERUP(tdi_STEPDOWNalgorithmCONTROL1p3_POWERUP_XU64),
.ten_STEPDOWNalgorithmCONTROL1p3_POWERUP(ten_STEPDOWNalgorithmCONTROL1p3_POWERUP_XU64)
);

dftprobe_XLOOP_XCONTROL_XU65 XU65 (
.i(net_312),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_FAULT(tdi_STEPDOWNalgorithmCONTROL1p3_FAULT_XU65),
.ten_STEPDOWNalgorithmCONTROL1p3_FAULT(ten_STEPDOWNalgorithmCONTROL1p3_FAULT_XU65)
);

dftprobe_XLOOP_XCONTROL_XU66 XU66 (
.i(net_311),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_READY(tdi_STEPDOWNalgorithmCONTROL1p3_READY_XU66),
.ten_STEPDOWNalgorithmCONTROL1p3_READY(ten_STEPDOWNalgorithmCONTROL1p3_READY_XU66)
);

dftprobe_XLOOP_XCONTROL_XU67 XU67 (
.i(net_322),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_IDLE(tdi_STEPDOWNalgorithmCONTROL1p3_IDLE_XU67),
.ten_STEPDOWNalgorithmCONTROL1p3_IDLE(ten_STEPDOWNalgorithmCONTROL1p3_IDLE_XU67)
);

dftprobe_XLOOP_XCONTROL_XU68 XU68 (
.i(net_325),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_UNDEF5(tdi_STEPDOWNalgorithmCONTROL1p3_UNDEF5_XU68),
.ten_STEPDOWNalgorithmCONTROL1p3_UNDEF5(ten_STEPDOWNalgorithmCONTROL1p3_UNDEF5_XU68)
);

dftprobe_XLOOP_XCONTROL_XU69 XU69 (
.i(net_331),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_BOTTOM(tdi_STEPDOWNalgorithmCONTROL1p3_BOTTOM_XU69),
.ten_STEPDOWNalgorithmCONTROL1p3_BOTTOM(ten_STEPDOWNalgorithmCONTROL1p3_BOTTOM_XU69)
);

dftprobe_XLOOP_XCONTROL_XU70 XU70 (
.i(net_300),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_TOP(tdi_STEPDOWNalgorithmCONTROL1p3_TOP_XU70),
.ten_STEPDOWNalgorithmCONTROL1p3_TOP(ten_STEPDOWNalgorithmCONTROL1p3_TOP_XU70)
);

dftprobe_XLOOP_XCONTROL_XU71 XU71 (
.i(topstate),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_topstate(tdi_STEPDOWNalgorithmCONTROL1p3_topstate_XU71),
.ten_STEPDOWNalgorithmCONTROL1p3_topstate(ten_STEPDOWNalgorithmCONTROL1p3_topstate_XU71)
);

dftprobe_XLOOP_XCONTROL_XU72 XU72 (
.i(botstate),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_botstate(tdi_STEPDOWNalgorithmCONTROL1p3_botstate_XU72),
.ten_STEPDOWNalgorithmCONTROL1p3_botstate(ten_STEPDOWNalgorithmCONTROL1p3_botstate_XU72)
);

dftprobe_XLOOP_XCONTROL_XU73 XU73 (
.i(fault_controller),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCONTROL1p3_fault_controller(tdi_STEPDOWNalgorithmCONTROL1p3_fault_controller_XU73),
.ten_STEPDOWNalgorithmCONTROL1p3_fault_controller(ten_STEPDOWNalgorithmCONTROL1p3_fault_controller_XU73)
);

DFTtm8d dft_hex0x2 (
.G(CELG59462),
.V(CELV96848),
.a({a1,a0}),
.SUB(CELSUB40948),
.tdi({tdi_STEPDOWNalgorithmCONTROL1p3_TOP_XU70,tdi_STEPDOWNalgorithmCONTROL1p3_BOTTOM_XU69,tdi_STEPDOWNalgorithmCONTROL1p3_UNDEF5_XU68,tdi_STEPDOWNalgorithmCONTROL1p3_IDLE_XU67,tdi_STEPDOWNalgorithmCONTROL1p3_READY_XU66,tdi_STEPDOWNalgorithmCONTROL1p3_FAULT_XU65,tdi_STEPDOWNalgorithmCONTROL1p3_POWERUP_XU64,tdi_STEPDOWNalgorithmCONTROL1p3_OFF_XU63}),
.tdo(tdo),
.ten({ten_STEPDOWNalgorithmCONTROL1p3_TOP_XU70,ten_STEPDOWNalgorithmCONTROL1p3_BOTTOM_XU69,ten_STEPDOWNalgorithmCONTROL1p3_UNDEF5_XU68,ten_STEPDOWNalgorithmCONTROL1p3_IDLE_XU67,ten_STEPDOWNalgorithmCONTROL1p3_READY_XU66,ten_STEPDOWNalgorithmCONTROL1p3_FAULT_XU65,ten_STEPDOWNalgorithmCONTROL1p3_POWERUP_XU64,ten_STEPDOWNalgorithmCONTROL1p3_OFF_XU63}),
.tma({a0,a0,a0,a0,a0,a0,a1,a0}),
.tmi(tmi[4:0])
);

DFTtm8d dft_hex0x3 (
.G(CELG59462),
.V(CELV96848),
.a({b1,b0}),
.SUB(CELSUB40948),
.tdi({b0,b0,b0,b0,b0,tdi_STEPDOWNalgorithmCONTROL1p3_fault_controller_XU73,tdi_STEPDOWNalgorithmCONTROL1p3_botstate_XU72,tdi_STEPDOWNalgorithmCONTROL1p3_topstate_XU71}),
.tdo(tdo),
.ten({noconn_dft_hex0x3_ten_7,noconn_dft_hex0x3_ten_6,noconn_dft_hex0x3_ten_5,noconn_dft_hex0x3_ten_4,noconn_dft_hex0x3_ten_3,ten_STEPDOWNalgorithmCONTROL1p3_fault_controller_XU73,ten_STEPDOWNalgorithmCONTROL1p3_botstate_XU72,ten_STEPDOWNalgorithmCONTROL1p3_topstate_XU71}),
.tma({b0,b0,b0,b0,b0,b0,b1,b1}),
.tmi(tmi[4:0])
);

STONEnoconn XNCnoconn_dft_hex0x3_ten_3 (
.noconn(noconn_dft_hex0x3_ten_3)
);

STONEnoconn XNCnoconn_dft_hex0x3_ten_4 (
.noconn(noconn_dft_hex0x3_ten_4)
);

STONEnoconn XNCnoconn_dft_hex0x3_ten_5 (
.noconn(noconn_dft_hex0x3_ten_5)
);

STONEnoconn XNCnoconn_dft_hex0x3_ten_6 (
.noconn(noconn_dft_hex0x3_ten_6)
);

STONEnoconn XNCnoconn_dft_hex0x3_ten_7 (
.noconn(noconn_dft_hex0x3_ten_7)
);

endmodule

