module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU37 (i,tdi_SOFTSTARTinternalNOFAULT_DONE,ten_SOFTSTARTinternalNOFAULT_DONE,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTinternalNOFAULT_DONE;
input  ten_SOFTSTARTinternalNOFAULT_DONE;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

