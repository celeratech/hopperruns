//Celera:currentmirror1_XLOOP_XREGULATION_XU2_XGMCURRENT
//Celera Confidential Symbol Generator
//Polarity: source, Maximum Current: 20, Number of outputs: 1, DFT: no, Max Vout: 6
//GAIN0:2.5, TYPE0:source
module currentmirror1_XLOOP_XREGULATION_XU2_XGMCURRENT (SIMPV,CELSUB,enable_currentmirror,ISET,ok_currentmirror,ten,
I0,
CELG);
input SIMPV;
input CELG;
input CELSUB;
input enable_currentmirror;
input ISET;
output ok_currentmirror;
input ten;
inout I0;
endmodule

