module dfthijack_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU9 (ENABLEpowergoodo,CELG,CELV,CELSUB,ten_ENABLEpowergoodenable,ten_ENABLEpowergoodstatus,ENABLEpowergood);
output  ENABLEpowergoodo;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_ENABLEpowergoodenable;
input  ten_ENABLEpowergoodstatus;
input  ENABLEpowergood;
endmodule

