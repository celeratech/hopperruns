//Celera:fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XTOPSW
//Celera Confidential Symbol Generator
//power NMOS:Ron:0.400 Ohm
//Vgs 6V Vds 30V
//Kelvin:no

module fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XTOPSW (GATE,SOURCE,DRAIN,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
endmodule

