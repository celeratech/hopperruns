//Celera:fet_fet_fetdriver_XLOOP_XDRIVER_XTOPDRIVER_XTSWDRIVER_Xpmos0_Xfet
//Celera Confidential Symbol Generator
//power PMOS:Ron:4.000 Ohm
//Vgs 6V Vds 6V
//Kelvin:no

module fet_fet_fetdriver_XLOOP_XDRIVER_XTOPDRIVER_XTSWDRIVER_Xpmos0_Xfet (GATE,SOURCE,DRAIN,PMOSiso6,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
input PMOSiso6;
endmodule

