module dftprobe_XLOOP_XREG_XDEBUG_XU8 (i,TAI_REGref,ten_REGref,CELG,CELSUB,CELV);
input  i;
output  TAI_REGref;
input  ten_REGref;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

