//Celera:nor2_XLOOP_XCONTROL_XU31_XU11
//Celera Confidential Symbol Generator
//nor2
module nor2_XLOOP_XCONTROL_XU31_XU11 (CELV,CELG,i0,i1,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input SUB;
output o;
endmodule

