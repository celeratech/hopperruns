module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU35 (i,tdi_SOFTSTARTinternalNOFAULT_OFF,ten_SOFTSTARTinternalNOFAULT_OFF,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTinternalNOFAULT_OFF;
input  ten_SOFTSTARTinternalNOFAULT_OFF;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

