//Celera:delayfixed_XLOOP_XCONTROL_XU55_XU7
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:both
module delayfixed_XLOOP_XCONTROL_XU55_XU7 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

