//Celera:timingskew_XLOOP_XDRIVER_XBOTSW_XU18
//Celera Confidential Symbol Generator
//TYPE:rise Bits:4 with 2.0ns LSB
module timingskew_XLOOP_XDRIVER_XBOTSW_XU18 (CELV,in,out,
factory_timingskew,
CELG,CELSUB);
input CELV;
input in;
output out;
input [3:0] factory_timingskew;
input CELG;
input CELSUB;
endmodule

