module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU82 (i,tdi_STEPDOWNalgorithmCORE0p0_RUN,ten_STEPDOWNalgorithmCORE0p0_RUN,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_RUN;
input  ten_STEPDOWNalgorithmCORE0p0_RUN;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

