module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU72 (i,tdi_STEPDOWNalgorithmCONTROL0p2_TOP,ten_STEPDOWNalgorithmCONTROL0p2_TOP,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_TOP;
input  ten_STEPDOWNalgorithmCONTROL0p2_TOP;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

