module dftprobe_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU13 (i,TAI_REGULATIONslope,ten_REGULATIONslope,CELG,CELSUB,CELV);
input  i;
output  TAI_REGULATIONslope;
input  ten_REGULATIONslope;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

