module dftprobe_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU3 (i,tdi_POWERGOODoutput,ten_POWERGOODoutput,CELG,CELSUB,CELV);
input  i;
output  tdi_POWERGOODoutput;
input  ten_POWERGOODoutput;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

