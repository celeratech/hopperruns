//Celera:timingskew_XLOOP_XDRIVER_XBOTDRIVER_XU41
//Celera Confidential Symbol Generator
//TYPE:fall Bits:5 with 8.0ns LSB
module timingskew_XLOOP_XDRIVER_XBOTDRIVER_XU41 (CELV,in,out,
factory_timingskew,
CELG,CELSUB);
input CELV;
input in;
output out;
input [4:0] factory_timingskew;
input CELG;
input CELSUB;
endmodule

