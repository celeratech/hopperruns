//Celera:currentgenerator_currentlimitfet_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWILIM_Xcg
//Celera Confidential Symbol Generator
//Number of outputs: 1, Max Vout: 6V, Accuracy: no%, Temperature Coefficient: zero, Temperature Gain: 3, DFT: no
//POLARITY0:source, OUTPUT0:2.83
module currentgenerator_currentlimitfet_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWILIM_Xcg (CELV,SUB,enable_currentgenerator,ten,IP,ok_currentgenerator,
I0,
CELG);
input CELV;
input CELG;
input SUB;
input enable_currentgenerator;
input IP;
output ok_currentgenerator;
input ten;
inout I0;
endmodule

