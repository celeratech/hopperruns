//Celera:inv_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU8_XU53
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU8_XU53 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

