module dftprobe_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU15 (i,tdi_botswipeak,ten_botswipeak,CELG,CELSUB,CELV);
input  i;
output  tdi_botswipeak;
input  ten_botswipeak;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

