// ------------------------ Module Definitions -----------
module nand3_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU5_XU4 (CELV,CELG,i0,i1,i2,o,SUB);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU5_XU5 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

// ------------------------ Module Verilog ---------------
module VESPAasmINPUT2_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU5 (o, i0, i1, Tstate, CELG59462, CELV96848, CELSUB40948);
output  o;
input  i0;
input  i1;
input  Tstate;
input  CELG59462;
input  CELV96848;
input  CELSUB40948;


// ------------------------ Wires ------------------------

// ------------------------ Networks ---------------------
nand3_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU5_XU4 XU4 (
.o(net_5),
.i0(Tstate),
.i1(i1),
.i2(i0),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU5_XU5 XU5 (
.i(net_5),
.o(o),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

endmodule

