//Celera:delay0_delayfixed_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU9_XU14_delay0
//TYPE: fixed 5ns
module delay0_delayfixed_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU9_XU14_delay0 (i, CELV, o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELSUB;
input CELG;
endmodule

