module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU77 (i,tdi_STEPDOWNalgorithmCONTROL0p2_topstate,ten_STEPDOWNalgorithmCONTROL0p2_topstate,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_topstate;
input  ten_STEPDOWNalgorithmCONTROL0p2_topstate;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

