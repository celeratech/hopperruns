//Celera:dbuf_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU8_XU55
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU8_XU55 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

