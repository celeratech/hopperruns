//Celera:switchideal_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU7
//Celera Confidential Symbol Generator
//1000 Ohm transmissionSwitch
module switchideal_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU7 (CELV,O,I,enable_switch,CELG,CELSUB);
input CELV;
input I;
input enable_switch;
inout O;
input CELG;
input CELSUB;
endmodule

