//Celera:bgcomp_XU1_XSERVICE_XBIASSERVICE_XU2
//Celera Confidential Symbol Generator
//Trip threshold: 1.5V, Maximum Supply Voltage: 30V, Maximum Input Voltage:30V
//Logic shift output:no, Trim trip threshold: yes, Enable pin: no, DFT: no
module bgcomp_XU1_XSERVICE_XBIASSERVICE_XU2 (CELSUB,CELPOS,IN,out,global_bgcomp,
trim_bgcomp,
CELG);
input CELSUB;
input CELPOS;
input IN;
output out;
input global_bgcomp;
input [7:0] trim_bgcomp;
input CELG;
endmodule

