module dftprobe_XLOOP_XDRIVER_XDEBUG_XU12 (i,tdi_DRVstartup,ten_DRVstartup,CELG,CELSUB,CELV);
input  i;
output  tdi_DRVstartup;
input  ten_DRVstartup;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

