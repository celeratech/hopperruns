//Celera:timingskew_XU1_XSTEPDOWN_XCORESTATE_XU32_XU35
//Celera Confidential Symbol Generator
//TYPE:rise Bits:2 with 2.0ns LSB
module timingskew_XU1_XSTEPDOWN_XCORESTATE_XU32_XU35 (CELV,in,out,
s,
CELG,CELSUB);
input CELV;
input in;
output out;
input [1:0] s;
input CELG;
input CELSUB;
endmodule

