//Celera:dbuf_XLOOP_XCONTROL_XU12_XU6
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XLOOP_XCONTROL_XU12_XU6 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

