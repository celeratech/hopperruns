module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU70 (i,tdi_STEPDOWNalgorithmCONTROL0p2_POWERUP,ten_STEPDOWNalgorithmCONTROL0p2_POWERUP,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_POWERUP;
input  ten_STEPDOWNalgorithmCONTROL0p2_POWERUP;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

