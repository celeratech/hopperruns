module dftprobe_XLOOP_XCONTROL_XU63 (i,tdi_STEPDOWNalgorithmCONTROL1p3_OFF,ten_STEPDOWNalgorithmCONTROL1p3_OFF,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_OFF;
input  ten_STEPDOWNalgorithmCONTROL1p3_OFF;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

