//Celera:padopendrain_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU14
//Celera Confidential Symbol Generator
//Open Drain output PAD with 6V, Ron 100 Ohms
//No Glitch filter
//ON Logic:noninvert polarity
//DFT:no TESTMODE:no RETURN PIN:no
module padopendrain_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU14 (CELV, input_padopendrain, PAD, 
CELG, SUB ); 
input CELV;
input input_padopendrain;
input CELG;
input SUB;
inout PAD;
endmodule

