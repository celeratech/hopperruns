module dftprobe_XU1_XSERVICE_XATESERVICE_XU12 (i,tdi_ok_service,ten_ok_service,CELG,CELSUB,CELV);
input  i;
output  tdi_ok_service;
input  ten_ok_service;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

