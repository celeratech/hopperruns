//Celera:pulsestretch_XU1_XSTEPDOWN_XFAULT_XU6_XU3
//Celera Confidential Symbol Generator
//VMAX:6PULSE STRETCH:10ns with 0ns delay
module pulsestretch_XU1_XSTEPDOWN_XFAULT_XU6_XU3 (CELV,in,out,porb,
CELG,CELSUB);
input CELV;
input in;
input porb;
output out;
input CELG;
input CELSUB;
endmodule

