//Celera:nand2_XU1_XSTEPDOWN_XLOOP_XFEEDBACK_XU2_XU18_XU52
//Celera Confidential Symbol Generator
//5V NAND2
module nand2_XU1_XSTEPDOWN_XLOOP_XFEEDBACK_XU2_XU18_XU52 (CELV,CELG,i0,i1,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input SUB;
output o;
endmodule

