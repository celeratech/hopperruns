// Celera Brick Generator Confidential
//CORE:singlepowerfetN
//NAME:fet_fet_XLOOP_XDRIVER_XTOPDRIVER_XTOPSWREP_Xfet
//GENERATOR REVISION:0.3.9
//FET TYPE:n
//ON RESISTANCE:0.100 Ohms
//VDS RATING:6V
//VGS RATING:6V
//BODY DIODE:yes
//DIODE DRIVE:diode
//REPLICA:no
//REPLICA GAIN:10
//KEVLIN:no
//DFT:no
//ROTATE:no

//Celera Confidential Do Not Copy NMOS
module an5g6dw1_124p4x0p2x6p0x1p0 (DRAIN,GATE,SOURCE,ISO,SUB);
input GATE;
input ISO;
input SUB;
inout SOURCE;
inout DRAIN;
endmodule

//Celera Confidential Do Not Copy fet_fet_XLOOP_XDRIVER_XTOPDRIVER_XTOPSWREP_Xfet
//Celera Confidential Symbol Generator
//power NMOS:Ron:0.100 Ohm
//Vgs 6V Vds 6V
//Kelvin:no

module fet_fet_XLOOP_XDRIVER_XTOPDRIVER_XTOPSWREP_Xfet (GATE,SOURCE,DRAIN,NMOSiso6,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
input NMOSiso6;

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos0(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos1(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos2(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos3(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos4(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos5(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos6(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos7(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos8(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos9(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos10(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos11(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos12(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos13(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos14(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos15(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos16(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos17(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos18(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos19(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos20(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos21(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos22(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos23(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos24(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos25(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos26(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos27(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos28(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos29(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos30(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos31(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos32(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos33(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos34(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos35(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos36(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos37(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos38(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos39(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos40(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos41(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos42(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos43(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos44(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos45(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos46(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos47(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos48(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos49(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos50(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos51(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos52(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy an5g6dw1_124p4x0p2x6p0x1p0
an5g6dw1_124p4x0p2x6p0x1p0 Xnmos53(
.DRAIN (DRAIN),
.GATE (GATE),
.SOURCE (SOURCE),
.ISO (NMOSiso6),
.SUB (SUB)
);
//,diesize,an5g6dw1_124p4x0p2x6p0x1p0

//Celera Confidential Do Not Copy Module End
//Celera Schematic Generator
endmodule
