module dftprobe_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU16 (i,tdi_REGULATIONgo,ten_REGULATIONgo,CELG,CELSUB,CELV);
input  i;
output  tdi_REGULATIONgo;
input  ten_REGULATIONgo;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

