//Celera:dbuf_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU11
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU11 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

