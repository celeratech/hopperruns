// ------------------------ Module Definitions -----------
module VESPAclockSYNC_XLOOP_XCONTROL_XU10 (din,out,clock,state,CELG59462,CELV96848,CELSUB40948);
  input  din;
  output  out;
  input  clock;
  input  state;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAclockSYNC_XLOOP_XCONTROL_XU11 (din,out,clock,state,CELG59462,CELV96848,CELSUB40948);
  input  din;
  output  out;
  input  clock;
  input  state;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSTATE8PS_XLOOP_XCONTROL_XU12 (r0,r1,r2,s0,s1,s2,porb,state0,state1,state2,state3,state4,state5,state6,state7,CELG59462,CELV96848,CELSUB40948);
  input  r0;
  input  r1;
  input  r2;
  input  s0;
  input  s1;
  input  s2;
  input  porb;
  output  state0;
  output  state1;
  output  state2;
  output  state3;
  output  state4;
  output  state5;
  output  state6;
  output  state7;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU13 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU15 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XLOOP_XCONTROL_XU17 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU20 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XLOOP_XCONTROL_XU22 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XLOOP_XCONTROL_XU25 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU28 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XLOOP_XCONTROL_XU30 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmPRIORITY3_XLOOP_XCONTROL_XU32 (i0,i1,i2,o0,o1,o2,Tstate,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  o0;
  output  o1;
  output  o2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmPRIORITY2_XLOOP_XCONTROL_XU33 (i0,i1,o0,o1,Tstate,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  o0;
  output  o1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmPRIORITY3_XLOOP_XCONTROL_XU34 (i0,i1,i2,o0,o1,o2,Tstate,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  o0;
  output  o1;
  output  o2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU35 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT4_XLOOP_XCONTROL_XU36 (o,i0,i1,i2,i3,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT2_XLOOP_XCONTROL_XU37 (o,i0,i1,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT2_XLOOP_XCONTROL_XU38 (o,i0,i1,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU39 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT3_XLOOP_XCONTROL_XU40 (o,i0,i1,i2,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT3_XLOOP_XCONTROL_XU41 (o,i0,i1,i2,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT3_XLOOP_XCONTROL_XU42 (o,i0,i1,i2,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT2_XLOOP_XCONTROL_XU43 (o,i0,i1,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU44 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU45 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU46 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XLOOP_XCONTROL_XU47 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR3_XLOOP_XCONTROL_XU48 (i0,i1,i2,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR2_XLOOP_XCONTROL_XU49 (i0,i1,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR5_XLOOP_XCONTROL_XU50 (i0,i1,i2,i3,i4,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR2_XLOOP_XCONTROL_XU51 (i0,i1,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR3_XLOOP_XCONTROL_XU52 (i0,i1,i2,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR3_XLOOP_XCONTROL_XU53 (i0,i1,i2,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_1_XLOOP_XCONTROL_XU54 (o,i0,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT2_1_XLOOP_XCONTROL_XU55 (o,i0,tstate0,tstate1,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  tstate0;
  input  tstate1;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_0_XLOOP_XCONTROL_XU56 (o,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAclocktree3_XLOOP_XCONTROL_XU8 (clock0,clock1,clock2,clocki,CELG59462,CELV96848,CELSUB40948);
  output  clock0;
  output  clock1;
  output  clock2;
  input  clocki;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAclockSYNC_XLOOP_XCONTROL_XU9 (din,out,clock,state,CELG59462,CELV96848,CELSUB40948);
  input  din;
  output  out;
  input  clock;
  input  state;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module inv_XLOOP_XCONTROL_XU1 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU2 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU3 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU4 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU5 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU6 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XLOOP_XCONTROL_XU7 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module delayfixed_XLOOP_XCONTROL_XU14 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU16 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU18 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU19 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU21 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU23 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU24 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU26 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU27 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU29 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XLOOP_XCONTROL_XU31 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

// ------------------------ Module Verilog ---------------
module STEPDOWNalgorithmCONTROL0p2_PYES_XLOOP_XCONTROL (porb, clock, botstate, topstate, CELG59462, CELV96848, go_driver, ok_driver, botswipeak, topswipeak, CELSUB40948, botswstatus, botswzcross, topswstatus, enable_driver, fault_control);
input  porb;
input  clock;
output  botstate;
output  topstate;
input  CELG59462;
input  CELV96848;
input  go_driver;
input  ok_driver;
input  botswipeak;
input  topswipeak;
input  CELSUB40948;
input  botswstatus;
input  botswzcross;
input  topswstatus;
input  enable_driver;
output  fault_control;


// ------------------------ Wires ------------------------

// ------------------------ Networks ---------------------
VESPAclockSYNC_XLOOP_XCONTROL_XU10 XU10 (
.din(net_289),
.out(net_290),
.clock(net_259),
.state(net_291),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAclockSYNC_XLOOP_XCONTROL_XU11 XU11 (
.din(net_305),
.out(net_306),
.clock(net_270),
.state(net_288),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSTATE8PS_XLOOP_XCONTROL_XU12 XU12 (
.r0(net_257),
.r1(net_281),
.r2(net_287),
.s0(net_260),
.s1(net_277),
.s2(net_283),
.porb(porb),
.state0(net_252),
.state1(net_261),
.state2(net_271),
.state3(net_258),
.state4(net_282),
.state5(net_284),
.state6(net_288),
.state7(net_291),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU13 XU13 (
.state(net_252),
.Tstate(net_262),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_273),
.tmin_delayoutput(net_272)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU15 XU15 (
.state(net_261),
.Tstate(net_292),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_293),
.tmin_delayoutput(net_294)
);

VESPAasmTIMERminmax_XLOOP_XCONTROL_XU17 XU17 (
.state(net_271),
.Tstate(net_300),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_307),
.t_delayinput(net_298),
.tmax_delayoutput(net_310),
.tmin_delayoutput(net_299)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU20 XU20 (
.state(net_258),
.Tstate(net_253),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_317),
.tmin_delayoutput(net_316)
);

VESPAasmTIMERminmax_XLOOP_XCONTROL_XU22 XU22 (
.state(net_282),
.Tstate(net_318),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_320),
.t_delayinput(net_322),
.tmax_delayoutput(net_321),
.tmin_delayoutput(net_319)
);

VESPAasmTIMERminmax_XLOOP_XCONTROL_XU25 XU25 (
.state(net_284),
.Tstate(net_327),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_330),
.t_delayinput(net_332),
.tmax_delayoutput(net_331),
.tmin_delayoutput(net_329)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU28 XU28 (
.state(net_288),
.Tstate(net_308),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_334),
.tmin_delayoutput(net_333)
);

VESPAasmTIMERminimum_XLOOP_XCONTROL_XU30 XU30 (
.state(net_291),
.Tstate(net_323),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_336),
.tmin_delayoutput(net_335)
);

VESPAasmPRIORITY3_XLOOP_XCONTROL_XU32 XU32 (
.i0(net_263),
.i1(net_274),
.i2(net_278),
.o0(net_264),
.o1(net_275),
.o2(net_279),
.Tstate(net_253),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmPRIORITY2_XLOOP_XCONTROL_XU33 XU33 (
.i0(net_306),
.i1(net_314),
.o0(net_311),
.o1(net_309),
.Tstate(net_308),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmPRIORITY3_XLOOP_XCONTROL_XU34 XU34 (
.i0(net_325),
.i1(net_326),
.i2(net_290),
.o0(net_256),
.o1(net_265),
.o2(net_324),
.Tstate(net_323),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU35 XU35 (
.o(net_255),
.i0(enable_driver),
.Tstate(net_262),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT4_XLOOP_XCONTROL_XU36 XU36 (
.o(net_250),
.i0(enable_driver),
.i1(ok_driver),
.i2(clock),
.i3(go_driver),
.Tstate(net_292),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT2_XLOOP_XCONTROL_XU37 XU37 (
.o(net_263),
.i0(topswipeak),
.i1(clock),
.Tstate(net_253),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT2_XLOOP_XCONTROL_XU38 XU38 (
.o(net_274),
.i0(net_269),
.i1(net_286),
.Tstate(net_253),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU39 XU39 (
.o(net_278),
.i0(net_296),
.Tstate(net_253),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT3_XLOOP_XCONTROL_XU40 XU40 (
.o(net_325),
.i0(botswzcross),
.i1(clock),
.i2(go_driver),
.Tstate(net_323),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT3_XLOOP_XCONTROL_XU41 XU41 (
.o(net_326),
.i0(net_304),
.i1(botswzcross),
.i2(net_296),
.Tstate(net_323),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT3_XLOOP_XCONTROL_XU42 XU42 (
.o(net_289),
.i0(net_304),
.i1(clock),
.i2(go_driver),
.Tstate(net_323),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT2_XLOOP_XCONTROL_XU43 XU43 (
.o(net_305),
.i0(go_driver),
.i1(clock),
.Tstate(net_308),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU44 XU44 (
.o(net_314),
.i0(net_315),
.Tstate(net_308),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU45 XU45 (
.o(net_312),
.i0(net_315),
.Tstate(net_300),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU46 XU46 (
.o(net_328),
.i0(net_320),
.Tstate(net_318),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XLOOP_XCONTROL_XU47 XU47 (
.o(net_276),
.i0(net_330),
.Tstate(net_327),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR3_XLOOP_XCONTROL_XU48 XU48 (
.i0(net_256),
.i1(net_265),
.i2(net_276),
.sr(net_257),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR2_XLOOP_XCONTROL_XU49 XU49 (
.i0(net_309),
.i1(net_312),
.sr(net_281),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR5_XLOOP_XCONTROL_XU50 XU50 (
.i0(net_324),
.i1(net_311),
.i2(net_309),
.i3(net_328),
.i4(net_276),
.sr(net_287),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR2_XLOOP_XCONTROL_XU51 XU51 (
.i0(net_255),
.i1(net_311),
.sr(net_260),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR3_XLOOP_XCONTROL_XU52 XU52 (
.i0(net_251),
.i1(net_328),
.i2(net_276),
.sr(net_277),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR3_XLOOP_XCONTROL_XU53 XU53 (
.i0(net_264),
.i1(net_275),
.i2(net_279),
.sr(net_283),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_1_XLOOP_XCONTROL_XU54 XU54 (
.o(topstate),
.i0(net_266),
.tstate(net_258),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT2_1_XLOOP_XCONTROL_XU55 XU55 (
.o(botstate),
.i0(net_302),
.tstate0(net_261),
.tstate1(net_291),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_0_XLOOP_XCONTROL_XU56 XU56 (
.o(fault_control),
.tstate(net_271),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAclocktree3_XLOOP_XCONTROL_XU8 XU8 (
.clock0(net_249),
.clock1(net_259),
.clock2(net_270),
.clocki(clock),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAclockSYNC_XLOOP_XCONTROL_XU9 XU9 (
.din(net_250),
.out(net_251),
.clock(net_249),
.state(net_261),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

inv_XLOOP_XCONTROL_XU1 XU1 (
.i(topswipeak),
.o(net_269),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU2 XU2 (
.i(clock),
.o(net_286),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU3 XU3 (
.i(go_driver),
.o(net_296),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU4 XU4 (
.i(botswipeak),
.o(net_304),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU5 XU5 (
.i(enable_driver),
.o(net_315),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU6 XU6 (
.i(botswstatus),
.o(net_266),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XLOOP_XCONTROL_XU7 XU7 (
.i(topswstatus),
.o(net_302),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

delayfixed_XLOOP_XCONTROL_XU14 XU14 (
.i(net_273),
.o(net_272),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU16 XU16 (
.i(net_293),
.o(net_294),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU18 XU18 (
.i(net_298),
.o(net_299),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU19 XU19 (
.i(net_298),
.o(net_310),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU21 XU21 (
.i(net_317),
.o(net_316),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU23 XU23 (
.i(net_322),
.o(net_319),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU24 XU24 (
.i(net_322),
.o(net_321),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU26 XU26 (
.i(net_332),
.o(net_329),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU27 XU27 (
.i(net_332),
.o(net_331),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU29 XU29 (
.i(net_334),
.o(net_333),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XLOOP_XCONTROL_XU31 XU31 (
.i(net_336),
.o(net_335),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

endmodule

