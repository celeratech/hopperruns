//Celera:tie_XLOOP_XCONTROL_XU31_XU8
//Celera Confidential Symbol Generator
//TIE
module tie_XLOOP_XCONTROL_XU31_XU8 (CELV,CELG,a0,SUB);
input CELV;
input CELG;
output a0;
input SUB;
endmodule

