//Celera Brick Generator Confidential
//CORE:resistordivider
//NAME:resistordivider_vbias_XU1_XSERVICE_XBIASSERVICE_XU1_XRuvlo
//GENERATOR REVISION:0.4.6
//VMAX:6V
//VTOP:6V
//TOTAL:6000.0
//DISCONNECT:no
//DISCONNECT TAP:top
//OUTPUTS:1
//TAP0:33.3%
//TAP1:99%
//TAP2:99%
//TAP3:99%
//TAP4:99%
//TAP5:99%
//TAP6:99%
//TAP7:99%

//Celera Confidential Do Not Copy STONEnoconn
//Verilog HDL for "Generate", "STONEnoconn" "functional"


module STONEnoconn ( noconn );

  input noconn;
endmodule

//Celera Confidential Do Not Copy Resistor Divider
module rlpp3000rpo8p8u1p0u (ISO,RP,RN);
input ISO;
inout RP;
inout RN;
endmodule

//Celera Confidential Do Not Copy resistordivider_vbias_XU1_XSERVICE_XBIASSERVICE_XU1_XRuvlo
//Celera Confidential Symbol Generator
//VMAX:6V R:6000.0KOhm 1Taps
module resistordivider_vbias_XU1_XSERVICE_XBIASSERVICE_XU1_XRuvlo (TOP,
TAP0,
CELG, BOTTOM);
inout TOP;
output TAP0;
input CELG;
inout BOTTOM;

//Celera Confidential Do Not Copy RTOP
rlpp3000rpo8p8u1p0u XRTOP_0(
.RP (TOP),
.RN (TOPTAP0_1),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_1(
.RP (TOPTAP0_1),
.RN (TOPTAP0_2),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_2(
.RP (TOPTAP0_2),
.RN (TOPTAP0_3),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_3(
.RP (TOPTAP0_3),
.RN (TOPTAP0_4),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_4(
.RP (TOPTAP0_4),
.RN (TOPTAP0_5),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_5(
.RP (TOPTAP0_5),
.RN (TOPTAP0_6),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_6(
.RP (TOPTAP0_6),
.RN (TOPTAP0_7),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_7(
.RP (TOPTAP0_7),
.RN (TOPTAP0_8),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_8(
.RP (TOPTAP0_8),
.RN (TOPTAP0_9),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_9(
.RP (TOPTAP0_9),
.RN (TOPTAP0_10),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_10(
.RP (TOPTAP0_10),
.RN (TOPTAP0_11),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_11(
.RP (TOPTAP0_11),
.RN (TOPTAP0_12),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_12(
.RP (TOPTAP0_12),
.RN (TOPTAP0_13),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_13(
.RP (TOPTAP0_13),
.RN (TOPTAP0_14),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_14(
.RP (TOPTAP0_14),
.RN (TOPTAP0_15),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_15(
.RP (TOPTAP0_15),
.RN (TOPTAP0_16),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_16(
.RP (TOPTAP0_16),
.RN (TOPTAP0_17),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_17(
.RP (TOPTAP0_17),
.RN (TOPTAP0_18),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_18(
.RP (TOPTAP0_18),
.RN (TOPTAP0_19),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_19(
.RP (TOPTAP0_19),
.RN (TOPTAP0_20),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_20(
.RP (TOPTAP0_20),
.RN (TOPTAP0_21),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_21(
.RP (TOPTAP0_21),
.RN (TOPTAP0_22),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_22(
.RP (TOPTAP0_22),
.RN (TOPTAP0_23),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_23(
.RP (TOPTAP0_23),
.RN (TOPTAP0_24),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_24(
.RP (TOPTAP0_24),
.RN (TOPTAP0_25),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_25(
.RP (TOPTAP0_25),
.RN (TOPTAP0_26),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_26(
.RP (TOPTAP0_26),
.RN (TOPTAP0_27),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_27(
.RP (TOPTAP0_27),
.RN (TOPTAP0_28),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_28(
.RP (TOPTAP0_28),
.RN (TOPTAP0_29),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_29(
.RP (TOPTAP0_29),
.RN (TOPTAP0_30),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_30(
.RP (TOPTAP0_30),
.RN (TOPTAP0_31),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_31(
.RP (TOPTAP0_31),
.RN (TOPTAP0_32),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_32(
.RP (TOPTAP0_32),
.RN (TOPTAP0_33),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_33(
.RP (TOPTAP0_33),
.RN (TOPTAP0_34),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_34(
.RP (TOPTAP0_34),
.RN (TOPTAP0_35),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_35(
.RP (TOPTAP0_35),
.RN (TOPTAP0_36),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_36(
.RP (TOPTAP0_36),
.RN (TOPTAP0_37),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_37(
.RP (TOPTAP0_37),
.RN (TOPTAP0_38),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_38(
.RP (TOPTAP0_38),
.RN (TOPTAP0_39),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_39(
.RP (TOPTAP0_39),
.RN (TOPTAP0_40),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_40(
.RP (TOPTAP0_40),
.RN (TOPTAP0_41),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_41(
.RP (TOPTAP0_41),
.RN (TOPTAP0_42),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_42(
.RP (TOPTAP0_42),
.RN (TOPTAP0_43),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_43(
.RP (TOPTAP0_43),
.RN (TOPTAP0_44),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_44(
.RP (TOPTAP0_44),
.RN (TOPTAP0_45),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_45(
.RP (TOPTAP0_45),
.RN (TOPTAP0_46),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_46(
.RP (TOPTAP0_46),
.RN (TOPTAP0_47),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_47(
.RP (TOPTAP0_47),
.RN (TOPTAP0_48),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_48(
.RP (TOPTAP0_48),
.RN (TOPTAP0_49),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_49(
.RP (TOPTAP0_49),
.RN (TOPTAP0_50),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_50(
.RP (TOPTAP0_50),
.RN (TOPTAP0_51),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_51(
.RP (TOPTAP0_51),
.RN (TOPTAP0_52),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_52(
.RP (TOPTAP0_52),
.RN (TOPTAP0_53),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_53(
.RP (TOPTAP0_53),
.RN (TOPTAP0_54),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_54(
.RP (TOPTAP0_54),
.RN (TOPTAP0_55),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_55(
.RP (TOPTAP0_55),
.RN (TOPTAP0_56),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_56(
.RP (TOPTAP0_56),
.RN (TOPTAP0_57),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_57(
.RP (TOPTAP0_57),
.RN (TOPTAP0_58),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_58(
.RP (TOPTAP0_58),
.RN (TOPTAP0_59),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_59(
.RP (TOPTAP0_59),
.RN (TOPTAP0_60),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_60(
.RP (TOPTAP0_60),
.RN (TOPTAP0_61),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_61(
.RP (TOPTAP0_61),
.RN (TOPTAP0_62),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_62(
.RP (TOPTAP0_62),
.RN (TOPTAP0_63),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_63(
.RP (TOPTAP0_63),
.RN (TOPTAP0_64),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_64(
.RP (TOPTAP0_64),
.RN (TOPTAP0_65),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_65(
.RP (TOPTAP0_65),
.RN (TOPTAP0_66),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_66(
.RP (TOPTAP0_66),
.RN (TOPTAP0_67),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_67(
.RP (TOPTAP0_67),
.RN (TOPTAP0_68),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_68(
.RP (TOPTAP0_68),
.RN (TOPTAP0_69),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_69(
.RP (TOPTAP0_69),
.RN (TOPTAP0_70),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_70(
.RP (TOPTAP0_70),
.RN (TOPTAP0_71),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_71(
.RP (TOPTAP0_71),
.RN (TOPTAP0_72),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_72(
.RP (TOPTAP0_72),
.RN (TOPTAP0_73),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_73(
.RP (TOPTAP0_73),
.RN (TOPTAP0_74),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_74(
.RP (TOPTAP0_74),
.RN (TOPTAP0_75),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_75(
.RP (TOPTAP0_75),
.RN (TOPTAP0_76),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_76(
.RP (TOPTAP0_76),
.RN (TOPTAP0_77),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_77(
.RP (TOPTAP0_77),
.RN (TOPTAP0_78),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_78(
.RP (TOPTAP0_78),
.RN (TOPTAP0_79),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_79(
.RP (TOPTAP0_79),
.RN (TOPTAP0_80),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_80(
.RP (TOPTAP0_80),
.RN (TOPTAP0_81),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_81(
.RP (TOPTAP0_81),
.RN (TOPTAP0_82),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_82(
.RP (TOPTAP0_82),
.RN (TOPTAP0_83),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_83(
.RP (TOPTAP0_83),
.RN (TOPTAP0_84),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_84(
.RP (TOPTAP0_84),
.RN (TOPTAP0_85),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_85(
.RP (TOPTAP0_85),
.RN (TOPTAP0_86),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_86(
.RP (TOPTAP0_86),
.RN (TOPTAP0_87),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_87(
.RP (TOPTAP0_87),
.RN (TOPTAP0_88),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_88(
.RP (TOPTAP0_88),
.RN (TOPTAP0_89),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_89(
.RP (TOPTAP0_89),
.RN (TOPTAP0_90),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_90(
.RP (TOPTAP0_90),
.RN (TOPTAP0_91),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_91(
.RP (TOPTAP0_91),
.RN (TOPTAP0_92),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_92(
.RP (TOPTAP0_92),
.RN (TOPTAP0_93),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_93(
.RP (TOPTAP0_93),
.RN (TOPTAP0_94),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_94(
.RP (TOPTAP0_94),
.RN (TOPTAP0_95),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_95(
.RP (TOPTAP0_95),
.RN (TOPTAP0_96),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_96(
.RP (TOPTAP0_96),
.RN (TOPTAP0_97),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_97(
.RP (TOPTAP0_97),
.RN (TOPTAP0_98),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_98(
.RP (TOPTAP0_98),
.RN (TOPTAP0_99),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_99(
.RP (TOPTAP0_99),
.RN (TOPTAP0_100),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_100(
.RP (TOPTAP0_100),
.RN (TOPTAP0_101),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_101(
.RP (TOPTAP0_101),
.RN (TOPTAP0_102),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_102(
.RP (TOPTAP0_102),
.RN (TOPTAP0_103),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_103(
.RP (TOPTAP0_103),
.RN (TOPTAP0_104),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_104(
.RP (TOPTAP0_104),
.RN (TOPTAP0_105),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_105(
.RP (TOPTAP0_105),
.RN (TOPTAP0_106),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_106(
.RP (TOPTAP0_106),
.RN (TOPTAP0_107),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_107(
.RP (TOPTAP0_107),
.RN (TOPTAP0_108),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_108(
.RP (TOPTAP0_108),
.RN (TOPTAP0_109),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_109(
.RP (TOPTAP0_109),
.RN (TOPTAP0_110),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_110(
.RP (TOPTAP0_110),
.RN (TOPTAP0_111),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_111(
.RP (TOPTAP0_111),
.RN (TOPTAP0_112),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_112(
.RP (TOPTAP0_112),
.RN (TOPTAP0_113),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_113(
.RP (TOPTAP0_113),
.RN (TOPTAP0_114),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_114(
.RP (TOPTAP0_114),
.RN (TOPTAP0_115),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_115(
.RP (TOPTAP0_115),
.RN (TOPTAP0_116),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_116(
.RP (TOPTAP0_116),
.RN (TOPTAP0_117),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_117(
.RP (TOPTAP0_117),
.RN (TOPTAP0_118),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_118(
.RP (TOPTAP0_118),
.RN (TOPTAP0_119),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_119(
.RP (TOPTAP0_119),
.RN (TOPTAP0_120),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_120(
.RP (TOPTAP0_120),
.RN (TOPTAP0_121),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_121(
.RP (TOPTAP0_121),
.RN (TOPTAP0_122),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_122(
.RP (TOPTAP0_122),
.RN (TOPTAP0_123),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_123(
.RP (TOPTAP0_123),
.RN (TOPTAP0_124),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_124(
.RP (TOPTAP0_124),
.RN (TOPTAP0_125),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_125(
.RP (TOPTAP0_125),
.RN (TOPTAP0_126),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_126(
.RP (TOPTAP0_126),
.RN (TOPTAP0_127),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_127(
.RP (TOPTAP0_127),
.RN (TOPTAP0_128),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTOP_128(
.RP (TOPTAP0_128),
.RN (TAP0),
.ISO (CELG)
);

//Celera Confidential Do Not Copy //DieSize,rlpp3000rpo8p8u1p0u

//Die Size Calculator rlpp3000rpo8p8u1p0u
//,diesize,rlpp3000rpo8p8u1p0u,129

//Celera Confidential Do Not Copy RTAP0
rlpp3000rpo8p8u1p0u XRTAP0_0(
.RP (TAP0),
.RN (TAP0BOTTOM_1),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_1(
.RP (TAP0BOTTOM_1),
.RN (TAP0BOTTOM_2),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_2(
.RP (TAP0BOTTOM_2),
.RN (TAP0BOTTOM_3),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_3(
.RP (TAP0BOTTOM_3),
.RN (TAP0BOTTOM_4),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_4(
.RP (TAP0BOTTOM_4),
.RN (TAP0BOTTOM_5),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_5(
.RP (TAP0BOTTOM_5),
.RN (TAP0BOTTOM_6),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_6(
.RP (TAP0BOTTOM_6),
.RN (TAP0BOTTOM_7),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_7(
.RP (TAP0BOTTOM_7),
.RN (TAP0BOTTOM_8),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_8(
.RP (TAP0BOTTOM_8),
.RN (TAP0BOTTOM_9),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_9(
.RP (TAP0BOTTOM_9),
.RN (TAP0BOTTOM_10),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_10(
.RP (TAP0BOTTOM_10),
.RN (TAP0BOTTOM_11),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_11(
.RP (TAP0BOTTOM_11),
.RN (TAP0BOTTOM_12),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_12(
.RP (TAP0BOTTOM_12),
.RN (TAP0BOTTOM_13),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_13(
.RP (TAP0BOTTOM_13),
.RN (TAP0BOTTOM_14),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_14(
.RP (TAP0BOTTOM_14),
.RN (TAP0BOTTOM_15),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_15(
.RP (TAP0BOTTOM_15),
.RN (TAP0BOTTOM_16),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_16(
.RP (TAP0BOTTOM_16),
.RN (TAP0BOTTOM_17),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_17(
.RP (TAP0BOTTOM_17),
.RN (TAP0BOTTOM_18),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_18(
.RP (TAP0BOTTOM_18),
.RN (TAP0BOTTOM_19),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_19(
.RP (TAP0BOTTOM_19),
.RN (TAP0BOTTOM_20),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_20(
.RP (TAP0BOTTOM_20),
.RN (TAP0BOTTOM_21),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_21(
.RP (TAP0BOTTOM_21),
.RN (TAP0BOTTOM_22),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_22(
.RP (TAP0BOTTOM_22),
.RN (TAP0BOTTOM_23),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_23(
.RP (TAP0BOTTOM_23),
.RN (TAP0BOTTOM_24),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_24(
.RP (TAP0BOTTOM_24),
.RN (TAP0BOTTOM_25),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_25(
.RP (TAP0BOTTOM_25),
.RN (TAP0BOTTOM_26),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_26(
.RP (TAP0BOTTOM_26),
.RN (TAP0BOTTOM_27),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_27(
.RP (TAP0BOTTOM_27),
.RN (TAP0BOTTOM_28),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_28(
.RP (TAP0BOTTOM_28),
.RN (TAP0BOTTOM_29),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_29(
.RP (TAP0BOTTOM_29),
.RN (TAP0BOTTOM_30),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_30(
.RP (TAP0BOTTOM_30),
.RN (TAP0BOTTOM_31),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_31(
.RP (TAP0BOTTOM_31),
.RN (TAP0BOTTOM_32),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_32(
.RP (TAP0BOTTOM_32),
.RN (TAP0BOTTOM_33),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_33(
.RP (TAP0BOTTOM_33),
.RN (TAP0BOTTOM_34),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_34(
.RP (TAP0BOTTOM_34),
.RN (TAP0BOTTOM_35),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_35(
.RP (TAP0BOTTOM_35),
.RN (TAP0BOTTOM_36),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_36(
.RP (TAP0BOTTOM_36),
.RN (TAP0BOTTOM_37),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_37(
.RP (TAP0BOTTOM_37),
.RN (TAP0BOTTOM_38),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_38(
.RP (TAP0BOTTOM_38),
.RN (TAP0BOTTOM_39),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_39(
.RP (TAP0BOTTOM_39),
.RN (TAP0BOTTOM_40),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_40(
.RP (TAP0BOTTOM_40),
.RN (TAP0BOTTOM_41),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_41(
.RP (TAP0BOTTOM_41),
.RN (TAP0BOTTOM_42),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_42(
.RP (TAP0BOTTOM_42),
.RN (TAP0BOTTOM_43),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_43(
.RP (TAP0BOTTOM_43),
.RN (TAP0BOTTOM_44),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_44(
.RP (TAP0BOTTOM_44),
.RN (TAP0BOTTOM_45),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_45(
.RP (TAP0BOTTOM_45),
.RN (TAP0BOTTOM_46),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_46(
.RP (TAP0BOTTOM_46),
.RN (TAP0BOTTOM_47),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_47(
.RP (TAP0BOTTOM_47),
.RN (TAP0BOTTOM_48),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_48(
.RP (TAP0BOTTOM_48),
.RN (TAP0BOTTOM_49),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_49(
.RP (TAP0BOTTOM_49),
.RN (TAP0BOTTOM_50),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_50(
.RP (TAP0BOTTOM_50),
.RN (TAP0BOTTOM_51),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_51(
.RP (TAP0BOTTOM_51),
.RN (TAP0BOTTOM_52),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_52(
.RP (TAP0BOTTOM_52),
.RN (TAP0BOTTOM_53),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_53(
.RP (TAP0BOTTOM_53),
.RN (TAP0BOTTOM_54),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_54(
.RP (TAP0BOTTOM_54),
.RN (TAP0BOTTOM_55),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_55(
.RP (TAP0BOTTOM_55),
.RN (TAP0BOTTOM_56),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_56(
.RP (TAP0BOTTOM_56),
.RN (TAP0BOTTOM_57),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_57(
.RP (TAP0BOTTOM_57),
.RN (TAP0BOTTOM_58),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_58(
.RP (TAP0BOTTOM_58),
.RN (TAP0BOTTOM_59),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_59(
.RP (TAP0BOTTOM_59),
.RN (TAP0BOTTOM_60),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_60(
.RP (TAP0BOTTOM_60),
.RN (TAP0BOTTOM_61),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_61(
.RP (TAP0BOTTOM_61),
.RN (TAP0BOTTOM_62),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_62(
.RP (TAP0BOTTOM_62),
.RN (TAP0BOTTOM_63),
.ISO (CELG)
);
rlpp3000rpo8p8u1p0u XRTAP0_63(
.RP (TAP0BOTTOM_63),
.RN (BOTTOM),
.ISO (CELG)
);

//Celera Confidential Do Not Copy //DieSize,rlpp3000rpo8p8u1p0u

//Die Size Calculator rlpp3000rpo8p8u1p0u
//,diesize,rlpp3000rpo8p8u1p0u,64

//Celera Confidential Do Not Copy Module End
//Celera Schematic Generator
endmodule
