//Celera:resistor_XLOOP_XREG_XFREQ_XRDCGAIN
//Celera Confidential Symbol Generator
//RESISTOR:5000KOhm TYPE:poly DFT:no
module resistor_XLOOP_XREG_XFREQ_XRDCGAIN (RP,
CELG,
RN);
inout RP;
inout RN;
input CELG;
endmodule

