//Celera:fet_padopendrain_XU1_XSTEPDOWN_XPOWERGOOD_XU10_XU2_Xnmos
//Celera Confidential Symbol Generator
//power NMOS:Ron:50.000 Ohm
//Vgs 6V Vds 6V
//Kelvin:no

module fet_padopendrain_XU1_XSTEPDOWN_XPOWERGOOD_XU10_XU2_Xnmos (GATE,SOURCE,DRAIN,NMOSiso6,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input NMOSiso6;
input SUB;
endmodule

