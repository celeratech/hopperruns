//Celera:feedbackdivider_XU1_XSTEPDOWN_XLOOP_XFEEDBACK_XU1_XU2
//Celera Confidential Symbol Generator
//Type: control, Feedback Voltage: 1V, Disconnect Pin: pin, P Offset: 0%, N Offset: 0%, Bias Current: 5, DFT: no
//VOUT0:1.2V, VOUT1: 1.5V, VOUT2: 2V, VOUT3: 2.5V, VOUT4: 2.8V, VOUT5: 3V, VOUT6: 3.3V, VOUT7: 5V
module feedbackdivider_XU1_XSTEPDOWN_XLOOP_XFEEDBACK_XU1_XU2 (CELV,SUB,SENSE_FEEDBACKDIVIDER,FEEDBACKDIVIDER_FB,ten,RTN,
pin1,pin2,pin3,
enable_feedbackdivider,
CELG);
input CELV;
input SUB;
input SENSE_FEEDBACKDIVIDER;
output FEEDBACKDIVIDER_FB;
input ten;
input RTN;
input pin1;
input pin2;
input pin3;
input enable_feedbackdivider;
input CELG;
endmodule

