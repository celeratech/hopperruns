module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU79 (i,tdi_STEPDOWNalgorithmCORE0p0_POWERUP,ten_STEPDOWNalgorithmCORE0p0_POWERUP,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_POWERUP;
input  ten_STEPDOWNalgorithmCORE0p0_POWERUP;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

