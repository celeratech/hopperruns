module dftprobe_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU2 (i,tdi_REGULATIONstartup,ten_REGULATIONstartup,CELG,CELSUB,CELV);
input  i;
output  tdi_REGULATIONstartup;
input  ten_REGULATIONstartup;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

