module dfthijack_XLOOP_XREG_XDEBUG_XU4 (HJregeno,CELG,CELV,CELSUB,ten_HJregenenable,ten_HJregenstatus,HJregen);
output  HJregeno;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJregenenable;
input  ten_HJregenstatus;
input  HJregen;
endmodule

