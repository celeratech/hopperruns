module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU85 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_feedback,ten_STEPDOWNalgorithmCORE0p0_enable_feedback,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_enable_feedback;
input  ten_STEPDOWNalgorithmCORE0p0_enable_feedback;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

