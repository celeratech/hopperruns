//Celera:resistordivider_XLOOP_XREG_XFREQ_XU9
//Celera Confidential Symbol Generator
//VMAX:6V R:1000.0KOhm 1Taps
module resistordivider_XLOOP_XREG_XFREQ_XU9 (TOP,
TAP0,
CELG, BOTTOM);
inout TOP;
output TAP0;
input CELG;
inout BOTTOM;
endmodule

