module dftprobe1_XLOOP_XDRIVER_XDEBUG_XU10 (i,tdi_DRVtopswipeak,ten_DRVtopswipeak,CELG,CELSUB,CELV);
input  i;
output  tdi_DRVtopswipeak;
input  ten_DRVtopswipeak;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

