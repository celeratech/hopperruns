module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU76 (i,tdi_STEPDOWNalgorithmCONTROL0p2_BOTTOM,ten_STEPDOWNalgorithmCONTROL0p2_BOTTOM,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_BOTTOM;
input  ten_STEPDOWNalgorithmCONTROL0p2_BOTTOM;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

