//Celera:switchideal_XLOOP_XREG_XDEBUG_XU10
//Celera Confidential Symbol Generator
//1000 Ohm tswitchSwitch
module switchideal_XLOOP_XREG_XDEBUG_XU10 (CELV,O,I,enable_switch,CELG,CELSUB);
input CELV;
input I;
input enable_switch;
inout O;
input CELG;
input CELSUB;
endmodule

