//Celera:dff_XLOOP_XDRIVER_XTOPDRIVER_XU27
//Celera Confidential Symbol Generator
//DFF latch
module dff_XLOOP_XDRIVER_XTOPDRIVER_XU27 (CELV,CELG,d,rb,ck,q,qb,SUB );
input CELV;
input CELG;
input d;
input rb;
input ck;
input SUB;
output q;
output qb;
endmodule

