//Celera:dff_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU27
//Celera Confidential Symbol Generator
//DFF latch
module dff_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU27 (CELV,CELG,d,rb,ck,q,qb,SUB );
input CELV;
input CELG;
input d;
input rb;
input ck;
input SUB;
output q;
output qb;
endmodule

