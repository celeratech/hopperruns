// ------------------------ Module Definitions -----------
module nor2_XU1_XSTEPDOWN_XCORESTATE_XU65_XU2 (CELV,CELG,i0,i1,o,SUB);
  output  o;
  input  i0;
  input  i1;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XCORESTATE_XU65_XU6 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module dbuf_XU1_XSTEPDOWN_XCORESTATE_XU65_XU25 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

// ------------------------ Module Verilog ---------------
module VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU65 (i0, i1, sr, CELG59462, CELV96848, CELSUB40948);
input  i0;
input  i1;
output  sr;
input  CELG59462;
input  CELV96848;
input  CELSUB40948;


// ------------------------ Wires ------------------------

// ------------------------ Networks ---------------------
nor2_XU1_XSTEPDOWN_XCORESTATE_XU65_XU2 XU2 (
.o(net_4),
.i0(i0),
.i1(i1),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XCORESTATE_XU65_XU6 XU6 (
.i(net_4),
.o(net_5),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

dbuf_XU1_XSTEPDOWN_XCORESTATE_XU65_XU25 XU25 (
.i(net_5),
.o(sr),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

endmodule

