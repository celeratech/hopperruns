module dfthijack_XLOOP_XATE_XU7 (HJgodrivero,CELG,CELV,CELSUB,ten_HJgodriverenable,ten_HJgodriverstatus,HJgodriver);
output  HJgodrivero;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJgodriverenable;
input  ten_HJgodriverstatus;
input  HJgodriver;
endmodule

