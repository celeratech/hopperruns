module dftprobe_XLOOP_XCONTROL_XU66 (i,tdi_STEPDOWNalgorithmCONTROL1p3_READY,ten_STEPDOWNalgorithmCONTROL1p3_READY,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_READY;
input  ten_STEPDOWNalgorithmCONTROL1p3_READY;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

