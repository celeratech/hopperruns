//Celera:levelshifter0L2H_XLOOP_XDRIVER_XTOPDRIVER_XU2
//Celera Confidential Symbol Generator
//Direction: low2high, Maximum high voltage:36V 
//Enable pin:no
module levelshifter0L2H_XLOOP_XDRIVER_XTOPDRIVER_XU2 (SIMPV,CELSUB,HVPOS,HVNEG,in,out,
CELG);
input SIMPV;
input CELG;
input CELSUB;
input HVPOS;
input HVNEG;
input in;
output out;
endmodule

