module dfthijack_XU1_XSERVICE_XATESERVICE_XU22 (hjencoreo,CELG,CELV,CELSUB,ten_hjencoreenable,ten_hjencorestatus,hjencore);
output  hjencoreo;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_hjencoreenable;
input  ten_hjencorestatus;
input  hjencore;
endmodule

