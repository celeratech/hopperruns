//Celera:logicshifter0L2H_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xenable
//Logic Level shifter with Enable
module logicshifter0L2H_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xenable (enable_logicshifter,
HVPOS,HVNEG,SIMPV,
in,
out,
CELG,CELSUB);
input HVPOS;
input HVNEG;
input SIMPV;
input in;
output out;
input enable_logicshifter;
input CELSUB;
input CELG;
endmodule

