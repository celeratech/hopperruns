// Celera Brick Generator Confidential
//CORE:capacitorfixed
//NAME:capacitorfixed_slopecomp_XLOOP_XREGULATION_XU2_XU9_Xslc
//GENERATOR REVISION:0.3.4
//VALUE:20.00Kohms
//Initial Voltage:1V
//TYPE:mim
//VMAX:6V
//DFT:no
//KELVIN:no

//Celera Confidential Do Not Copy mim34_2f30p0x29p7
//Celera Confidential Symbol Generator
//Type mim :20.00pF Capacitor
module mim34_2f30p0x29p7 (CP, CN);
inout CP;
inout CN;
endmodule

//Celera Confidential Do Not Copy capacitorfixed_slopecomp_XLOOP_XREGULATION_XU2_XU9_Xslc
//Celera Confidential Symbol Generator
//CAPACITOR CONTROL:capacitor
//VALUE: 20.00pF TYPE:mim
module capacitorfixed_slopecomp_XLOOP_XREGULATION_XU2_XU9_Xslc (CP,
CN);
inout CP;
inout CN;

//Celera Confidential Do Not Copy Core_
mim34_2f30p0x29p7 XCore_0(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_1(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_2(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_3(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_4(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_5(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_6(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_7(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_8(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_9(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x29p7 XCore_10(
.CP (CP),
.CN (CN)
);

//Celera Confidential Do Not Copy //DieSize,mim34_2f30p0x29p7

//Die Size Calculator mim34_2f30p0x29p7
//,diesize,mim34_2f30p0x29p7,11

//Celera Confidential Do Not Copy Module End
//Celera Schematic Generator
endmodule
