module dftprobe_XU1_XSERVICE_XATESERVICE_XU3 (i,tdi_envbias,ten_envbias,CELG,CELSUB,CELV);
input  i;
output  tdi_envbias;
input  ten_envbias;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

