//Celera:inv_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU5_XU5
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSTEPDOWN_XPOWERGOOD_XU7_XU5_XU5 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

