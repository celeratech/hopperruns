//Celera:oneshot_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU9_XU13
//Celera Confidential Symbol Generator
//One Shot100ns OneShot - Bad Designer!!
module oneshot_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU9_XU13 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

