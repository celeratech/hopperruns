//Celera:inv_XLOOP_XREG_XFREQ_XU12
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XLOOP_XREG_XFREQ_XU12 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

