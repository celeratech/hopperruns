//Celera:dbuf_XLOOP_XREGULATION_XU2_XU10
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XLOOP_XREGULATION_XU2_XU10 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

