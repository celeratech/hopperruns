module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU77 (i,tdi_STEPDOWNalgorithmCORE0p0_DISCHARGE,ten_STEPDOWNalgorithmCORE0p0_DISCHARGE,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_DISCHARGE;
input  ten_STEPDOWNalgorithmCORE0p0_DISCHARGE;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

