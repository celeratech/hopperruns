//Celera:dbuf_XU1_XSTEPDOWN_XSOFTSTART_XU7_XU10_XU55
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XSOFTSTART_XU7_XU10_XU55 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

