//Celera:tie_XLOOP_XDRIVER_XBOTDRIVER_XU39
//Celera Confidential Symbol Generator
//TIE
module tie_XLOOP_XDRIVER_XBOTDRIVER_XU39 (CELV,CELG,a1,SUB);
input CELV;
input CELG;
output a1;
input SUB;
endmodule

