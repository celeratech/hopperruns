module dftprobe_XLOOP_XCONTROL_XU64 (i,tdi_STEPDOWNalgorithmCONTROL1p3_POWERUP,ten_STEPDOWNalgorithmCONTROL1p3_POWERUP,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_POWERUP;
input  ten_STEPDOWNalgorithmCONTROL1p3_POWERUP;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

