//Celera:delay0_delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU27_delay0
//TYPE: fixed 100ns
module delay0_delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU4_XU27_delay0 (i, CELV, o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELSUB;
input CELG;
endmodule

