module dftprobe_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU14 (i,TAI_REGULATIONref,ten_REGULATIONref,CELG,CELSUB,CELV);
input  i;
output  TAI_REGULATIONref;
input  ten_REGULATIONref;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

