module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU71 (i,tdi_STEPDOWNalgorithmCONTROL0p2_FAULT,ten_STEPDOWNalgorithmCONTROL0p2_FAULT,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_FAULT;
input  ten_STEPDOWNalgorithmCONTROL0p2_FAULT;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

