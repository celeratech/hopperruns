//Celera:dbuf_XU1_XSERVICE_XATESERVICE_XU9_XU55
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSERVICE_XATESERVICE_XU9_XU55 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

