//Celera:resistor_XLOOP_XREGULATION_XU2_XRZCOMP
//Celera Confidential Symbol Generator
//RESISTOR:200.00KOhm TYPE:poly Adjust:200.00Kohm DFT:no
module resistor_XLOOP_XREGULATION_XU2_XRZCOMP (RP,
CELV,
CELG,
CELSUB,
factory_adjust_resistor,
RN);
inout RP;
inout RN;
input CELV;
input CELG;
input CELSUB;
input [2:0] factory_adjust_resistor;
endmodule

