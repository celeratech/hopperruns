// ------------------------ Module Definitions -----------
module VESPAasmOUTPUT2_0_XU1_XSTEPDOWN_XCORESTATE_XU10 (o,tstate0,tstate1,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate0;
  input  tstate1;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmTIMERminimum_XU1_XSTEPDOWN_XCORESTATE_XU11 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU13 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XU1_XSTEPDOWN_XCORESTATE_XU16 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU18 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU21 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU24 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminimum_XU1_XSTEPDOWN_XCORESTATE_XU27 (state,Tstate,CELG59462,CELV96848,CELSUB40948,tmin_delayinput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  tmin_delayinput;
  input  tmin_delayoutput;
endmodule

module VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU29 (state,Tstate,CELG59462,CELV96848,CELSUB40948,STATEtimeout,t_delayinput,tmax_delayoutput,tmin_delayoutput);
  input  state;
  output  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  output  STATEtimeout;
  output  t_delayinput;
  input  tmax_delayoutput;
  input  tmin_delayoutput;
endmodule

module VESPAasmPRIORITYD3_XU1_XSTEPDOWN_XCORESTATE_XU32 (i0,i1,i2,o0,o1,o2,Tstate,CELG59462,CELV96848,CELSUB40948,Tpriority0_0,Tpriority0_1,TpriorityX_0,TpriorityX_1,TpriorityX_2,TpriorityX_3);
  input  i0;
  input  i1;
  input  i2;
  output  o0;
  output  o1;
  output  o2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  input  Tpriority0_0;
  input  Tpriority0_1;
  input  TpriorityX_0;
  input  TpriorityX_1;
  input  TpriorityX_2;
  input  TpriorityX_3;
endmodule

module VESPAasmPRIORITYD2_XU1_XSTEPDOWN_XCORESTATE_XU35 (i0,i1,o0,o1,Tstate,CELG59462,CELV96848,CELSUB40948,Tpriority0_0,Tpriority0_1,TpriorityX_0,TpriorityX_1);
  input  i0;
  input  i1;
  output  o0;
  output  o1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  input  Tpriority0_0;
  input  Tpriority0_1;
  input  TpriorityX_0;
  input  TpriorityX_1;
endmodule

module VESPAasmPRIORITYD6_XU1_XSTEPDOWN_XCORESTATE_XU38 (i0,i1,i2,i3,i4,i5,o0,o1,o2,o3,o4,o5,Tstate,CELG59462,CELV96848,CELSUB40948,Tpriority0_0,Tpriority0_1,TpriorityX_0,TpriorityX_1,TpriorityX_2,TpriorityX_3,TpriorityX_4,TpriorityX_5,TpriorityX_6,TpriorityX_7,TpriorityY_0,TpriorityY_1);
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  input  i5;
  output  o0;
  output  o1;
  output  o2;
  output  o3;
  output  o4;
  output  o5;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  input  Tpriority0_0;
  input  Tpriority0_1;
  input  TpriorityX_0;
  input  TpriorityX_1;
  input  TpriorityX_2;
  input  TpriorityX_3;
  input  TpriorityX_4;
  input  TpriorityX_5;
  input  TpriorityX_6;
  input  TpriorityX_7;
  input  TpriorityY_0;
  input  TpriorityY_1;
endmodule

module VESPAasmPRIORITYD2_XU1_XSTEPDOWN_XCORESTATE_XU42 (i0,i1,o0,o1,Tstate,CELG59462,CELV96848,CELSUB40948,Tpriority0_0,Tpriority0_1,TpriorityX_0,TpriorityX_1);
  input  i0;
  input  i1;
  output  o0;
  output  o1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
  input  Tpriority0_0;
  input  Tpriority0_1;
  input  TpriorityX_0;
  input  TpriorityX_1;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU45 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT2_XU1_XSTEPDOWN_XCORESTATE_XU46 (o,i0,i1,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU47 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT3_XU1_XSTEPDOWN_XCORESTATE_XU48 (o,i0,i1,i2,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT4_XU1_XSTEPDOWN_XCORESTATE_XU49 (o,i0,i1,i2,i3,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU50 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT5_XU1_XSTEPDOWN_XCORESTATE_XU51 (o,i0,i1,i2,i3,i4,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU52 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU53 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU54 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU55 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU56 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU57 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU58 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU59 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU60 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU61 (o,i0,Tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  Tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR6_XU1_XSTEPDOWN_XCORESTATE_XU62 (i0,i1,i2,i3,i4,i5,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  input  i5;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR9_XU1_XSTEPDOWN_XCORESTATE_XU63 (i0,i1,i2,i3,i4,i5,i6,i7,i8,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  input  i2;
  input  i3;
  input  i4;
  input  i5;
  input  i6;
  input  i7;
  input  i8;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU64 (i0,i1,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU65 (i0,i1,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU66 (i0,i1,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU67 (i0,i1,sr,CELG59462,CELV96848,CELSUB40948);
  input  i0;
  input  i1;
  output  sr;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT3_0_XU1_XSTEPDOWN_XCORESTATE_XU68 (o,tstate0,tstate1,tstate2,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate0;
  input  tstate1;
  input  tstate2;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT2_0_XU1_XSTEPDOWN_XCORESTATE_XU69 (o,tstate0,tstate1,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate0;
  input  tstate1;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmSTATE8DF_XU1_XSTEPDOWN_XCORESTATE_XU7 (r0,r1,r2,s0,s1,s2,porb,state0,state1,state2,state3,state4,state5,state6,state7,CELG59462,CELV96848,hjconfig_0,hjconfig_1,hjconfig_2,hjconfig_3,CELSUB40948);
  input  r0;
  input  r1;
  input  r2;
  input  s0;
  input  s1;
  input  s2;
  input  porb;
  output  state0;
  output  state1;
  output  state2;
  output  state3;
  output  state4;
  output  state5;
  output  state6;
  output  state7;
  input  CELG59462;
  input  CELV96848;
  input  hjconfig_0;
  input  hjconfig_1;
  input  hjconfig_2;
  input  hjconfig_3;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_1_XU1_XSTEPDOWN_XCORESTATE_XU71 (o,i0,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  i0;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XCORESTATE_XU72 (o,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT3_0_XU1_XSTEPDOWN_XCORESTATE_XU74 (o,tstate0,tstate1,tstate2,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate0;
  input  tstate1;
  input  tstate2;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XCORESTATE_XU75 (o,tstate,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module VESPAasmOUTPUT5_0_XU1_XSTEPDOWN_XCORESTATE_XU9 (o,tstate0,tstate1,tstate2,tstate3,tstate4,CELG59462,CELV96848,CELSUB40948);
  output  o;
  input  tstate0;
  input  tstate1;
  input  tstate2;
  input  tstate3;
  input  tstate4;
  input  CELG59462;
  input  CELV96848;
  input  CELSUB40948;
endmodule

module inv_XU1_XSTEPDOWN_XCORESTATE_XU1 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XCORESTATE_XU2 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XCORESTATE_XU3 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XCORESTATE_XU4 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XCORESTATE_XU5 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XCORESTATE_XU6 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU12 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU14 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU15 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU17 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU19 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU20 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU22 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU23 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU25 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU26 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU28 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU30 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU31 (CELV,i,o,CELG,CELSUB);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU76 (i,tdi_STEPDOWNalgorithmCORE0p0_OFF,ten_STEPDOWNalgorithmCORE0p0_OFF,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_OFF;
  input  ten_STEPDOWNalgorithmCORE0p0_OFF;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU77 (i,tdi_STEPDOWNalgorithmCORE0p0_DISCHARGE,ten_STEPDOWNalgorithmCORE0p0_DISCHARGE,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_DISCHARGE;
  input  ten_STEPDOWNalgorithmCORE0p0_DISCHARGE;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU78 (i,tdi_STEPDOWNalgorithmCORE0p0_FAULT,ten_STEPDOWNalgorithmCORE0p0_FAULT,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_FAULT;
  input  ten_STEPDOWNalgorithmCORE0p0_FAULT;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU79 (i,tdi_STEPDOWNalgorithmCORE0p0_POWERUP,ten_STEPDOWNalgorithmCORE0p0_POWERUP,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_POWERUP;
  input  ten_STEPDOWNalgorithmCORE0p0_POWERUP;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU80 (i,tdi_STEPDOWNalgorithmCORE0p0_POWERDOWN,ten_STEPDOWNalgorithmCORE0p0_POWERDOWN,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_POWERDOWN;
  input  ten_STEPDOWNalgorithmCORE0p0_POWERDOWN;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU81 (i,tdi_STEPDOWNalgorithmCORE0p0_UNDEF5,ten_STEPDOWNalgorithmCORE0p0_UNDEF5,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_UNDEF5;
  input  ten_STEPDOWNalgorithmCORE0p0_UNDEF5;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU82 (i,tdi_STEPDOWNalgorithmCORE0p0_RUN,ten_STEPDOWNalgorithmCORE0p0_RUN,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_RUN;
  input  ten_STEPDOWNalgorithmCORE0p0_RUN;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU83 (i,tdi_STEPDOWNalgorithmCORE0p0_SOFTSTART,ten_STEPDOWNalgorithmCORE0p0_SOFTSTART,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_SOFTSTART;
  input  ten_STEPDOWNalgorithmCORE0p0_SOFTSTART;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU84 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_fault,ten_STEPDOWNalgorithmCORE0p0_enable_fault,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_enable_fault;
  input  ten_STEPDOWNalgorithmCORE0p0_enable_fault;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU85 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_feedback,ten_STEPDOWNalgorithmCORE0p0_enable_feedback,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_enable_feedback;
  input  ten_STEPDOWNalgorithmCORE0p0_enable_feedback;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU86 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_powergood,ten_STEPDOWNalgorithmCORE0p0_enable_powergood,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_enable_powergood;
  input  ten_STEPDOWNalgorithmCORE0p0_enable_powergood;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU87 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_softstart,ten_STEPDOWNalgorithmCORE0p0_enable_softstart,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_enable_softstart;
  input  ten_STEPDOWNalgorithmCORE0p0_enable_softstart;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU88 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_discharge,ten_STEPDOWNalgorithmCORE0p0_enable_discharge,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_enable_discharge;
  input  ten_STEPDOWNalgorithmCORE0p0_enable_discharge;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU89 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_regulation,ten_STEPDOWNalgorithmCORE0p0_enable_regulation,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_enable_regulation;
  input  ten_STEPDOWNalgorithmCORE0p0_enable_regulation;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU90 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_driver,ten_STEPDOWNalgorithmCORE0p0_enable_driver,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_enable_driver;
  input  ten_STEPDOWNalgorithmCORE0p0_enable_driver;
endmodule

module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU91 (i,tdi_STEPDOWNalgorithmCORE0p0_fault_core,ten_STEPDOWNalgorithmCORE0p0_fault_core,CELG,CELSUB,CELV);
  input  i;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_STEPDOWNalgorithmCORE0p0_fault_core;
  input  ten_STEPDOWNalgorithmCORE0p0_fault_core;
endmodule

//Verilog HDL for "DFT", "DFTtm8d" "functional"


module DFTtm8d ( a, ten, tdo, tmi, G, SUB, V, tdi, tma );

  input V;
  input  [7:0] tma;
  output  [7:0] ten;
  output  [1:0] a;
  inout tdo;
  input  [7:0] tdi;
  input G;
  input SUB;
  inout  [4:0] tmi;
endmodule


//Verilog HDL for "DRM", "drm32" "functional"


module drm32 ( V, G, SUB, tmi, bypload, lastdrm, id, por0, por1, por2, por3,
drm0, drm1, drm2, drm3, d1, d0 );

  input lastdrm;
  input V;
  output d1;
  input  [7:0] por3;
  output  [7:0] drm3;
  input  [7:0] id;
  output d0;
  output  [7:0] drm2;
  input  [7:0] por2;
  input  [7:0] por1;
  input bypload;
  output  [7:0] drm0;
  input  [7:0] por0;
  input G;
  output  [7:0] drm1;
  inout  [4:0] tmi;
  input SUB;
endmodule


//Verilog HDL for "Generate", "STONEnoconn" "functional"


module STONEnoconn ( noconn );

  input noconn;
endmodule


// ------------------------ Module Verilog ---------------
module STEPDOWNalgorithmCORE0p0_DYES_XU1_XSTEPDOWN_XCORESTATE (tdo, tmi, porb, ok_fault, CELG59462, CELV96848, ok_driver, fault_core, ok_service, CELSUB40948, ok_feedback, short_fault, enable_fault, ok_powergood, enable_driver, ok_regulation, done_discharge, done_softstart, enable_feedback, enable_discharge, enable_powergood, enable_softstart, enable_regulation);
inout  tdo;
inout [4:0] tmi;
input  porb;
input  ok_fault;
input  CELG59462;
input  CELV96848;
input  ok_driver;
output  fault_core;
input  ok_service;
input  CELSUB40948;
input  ok_feedback;
input  short_fault;
output  enable_fault;
input  ok_powergood;
output  enable_driver;
input  ok_regulation;
input  done_discharge;
input  done_softstart;
output  enable_feedback;
output  enable_discharge;
output  enable_powergood;
output  enable_softstart;
output  enable_regulation;


// ------------------------ Wires ------------------------
wire [4:0] tmi;
wire [1:0] a;
wire [7:0] tdi;
wire [7:0] ten;
wire [7:0] tma;
wire [7:0] id;
wire [7:0] drm0;
wire [7:0] drm1;
wire [7:0] drm2;
wire [7:0] drm3;
wire [7:0] por0;
wire [7:0] por1;
wire [7:0] por2;
wire [7:0] por3;

// ------------------------ Networks ---------------------
VESPAasmOUTPUT2_0_XU1_XSTEPDOWN_XCORESTATE_XU10 XU10 (
.o(enable_regulation),
.tstate0(net_394),
.tstate1(net_405),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmTIMERminimum_XU1_XSTEPDOWN_XCORESTATE_XU11 XU11 (
.state(net_385),
.Tstate(net_392),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_402),
.tmin_delayoutput(net_401)
);

VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU13 XU13 (
.state(net_391),
.Tstate(net_403),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_428),
.t_delayinput(net_424),
.tmax_delayoutput(net_429),
.tmin_delayoutput(net_425)
);

VESPAasmTIMERminimum_XU1_XSTEPDOWN_XCORESTATE_XU16 XU16 (
.state(net_400),
.Tstate(net_435),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_441),
.tmin_delayoutput(net_440)
);

VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU18 XU18 (
.state(net_390),
.Tstate(net_442),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_452),
.t_delayinput(net_455),
.tmax_delayoutput(net_454),
.tmin_delayoutput(net_451)
);

VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU21 XU21 (
.state(net_411),
.Tstate(net_458),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_460),
.t_delayinput(net_462),
.tmax_delayoutput(net_461),
.tmin_delayoutput(net_459)
);

VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU24 XU24 (
.state(net_415),
.Tstate(net_464),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_467),
.t_delayinput(net_470),
.tmax_delayoutput(net_469),
.tmin_delayoutput(net_466)
);

VESPAasmTIMERminimum_XU1_XSTEPDOWN_XCORESTATE_XU27 XU27 (
.state(net_394),
.Tstate(net_465),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.tmin_delayinput(net_477),
.tmin_delayoutput(net_476)
);

VESPAasmTIMERminmax_XU1_XSTEPDOWN_XCORESTATE_XU29 XU29 (
.state(net_405),
.Tstate(net_478),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.STATEtimeout(net_480),
.t_delayinput(net_482),
.tmax_delayoutput(net_481),
.tmin_delayoutput(net_479)
);

VESPAasmPRIORITYD3_XU1_XSTEPDOWN_XCORESTATE_XU32 XU32 (
.i0(net_406),
.i1(net_412),
.i2(net_416),
.o0(net_388),
.o1(net_393),
.o2(net_417),
.Tstate(net_403),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.Tpriority0_0(net_303),
.Tpriority0_1(net_304),
.TpriorityX_0(net_305),
.TpriorityX_1(net_306),
.TpriorityX_2(net_307),
.TpriorityX_3(net_308)
);

VESPAasmPRIORITYD2_XU1_XSTEPDOWN_XCORESTATE_XU35 XU35 (
.i0(net_444),
.i1(net_448),
.o0(net_445),
.o1(net_404),
.Tstate(net_442),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.Tpriority0_0(net_319),
.Tpriority0_1(net_320),
.TpriorityX_0(net_321),
.TpriorityX_1(net_322)
);

VESPAasmPRIORITYD6_XU1_XSTEPDOWN_XCORESTATE_XU38 XU38 (
.i0(net_468),
.i1(net_471),
.i2(net_472),
.i3(net_473),
.i4(net_474),
.i5(net_475),
.o0(net_443),
.o1(net_446),
.o2(net_449),
.o3(net_450),
.o4(net_453),
.o5(net_456),
.Tstate(net_465),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.Tpriority0_0(net_335),
.Tpriority0_1(net_336),
.TpriorityX_0(net_343),
.TpriorityX_1(net_344),
.TpriorityX_2(net_345),
.TpriorityX_3(net_346),
.TpriorityX_4(net_347),
.TpriorityX_5(net_348),
.TpriorityX_6(net_349),
.TpriorityX_7(net_350),
.TpriorityY_0(net_351),
.TpriorityY_1(net_352)
);

VESPAasmPRIORITYD2_XU1_XSTEPDOWN_XCORESTATE_XU42 XU42 (
.i0(net_483),
.i1(net_484),
.o0(net_407),
.o1(net_413),
.Tstate(net_478),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948),
.Tpriority0_0(net_359),
.Tpriority0_1(net_360),
.TpriorityX_0(net_367),
.TpriorityX_1(net_368)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU45 XU45 (
.o(net_387),
.i0(ok_service),
.Tstate(net_392),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT2_XU1_XSTEPDOWN_XCORESTATE_XU46 XU46 (
.o(net_406),
.i0(done_discharge),
.i1(net_436),
.Tstate(net_403),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU47 XU47 (
.o(net_412),
.i0(net_428),
.Tstate(net_403),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT3_XU1_XSTEPDOWN_XCORESTATE_XU48 XU48 (
.o(net_416),
.i0(done_discharge),
.i1(ok_feedback),
.i2(ok_service),
.Tstate(net_403),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT4_XU1_XSTEPDOWN_XCORESTATE_XU49 XU49 (
.o(net_444),
.i0(ok_feedback),
.i1(ok_driver),
.i2(ok_fault),
.i3(ok_service),
.Tstate(net_442),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU50 XU50 (
.o(net_448),
.i0(net_452),
.Tstate(net_442),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT5_XU1_XSTEPDOWN_XCORESTATE_XU51 XU51 (
.o(net_483),
.i0(done_softstart),
.i1(ok_feedback),
.i2(ok_driver),
.i3(ok_fault),
.i4(ok_service),
.Tstate(net_478),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU52 XU52 (
.o(net_484),
.i0(net_480),
.Tstate(net_478),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU53 XU53 (
.o(net_468),
.i0(short_fault),
.Tstate(net_465),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU54 XU54 (
.o(net_471),
.i0(net_398),
.Tstate(net_465),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU55 XU55 (
.o(net_472),
.i0(net_421),
.Tstate(net_465),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU56 XU56 (
.o(net_473),
.i0(net_432),
.Tstate(net_465),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU57 XU57 (
.o(net_474),
.i0(net_439),
.Tstate(net_465),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU58 XU58 (
.o(net_475),
.i0(net_447),
.Tstate(net_465),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU59 XU59 (
.o(net_457),
.i0(net_436),
.Tstate(net_435),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU60 XU60 (
.o(net_418),
.i0(net_467),
.Tstate(net_464),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmINPUT1_XU1_XSTEPDOWN_XCORESTATE_XU61 XU61 (
.o(net_463),
.i0(net_460),
.Tstate(net_458),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR6_XU1_XSTEPDOWN_XCORESTATE_XU62 XU62 (
.i0(net_388),
.i1(net_393),
.i2(net_404),
.i3(net_407),
.i4(net_413),
.i5(net_418),
.sr(net_389),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR9_XU1_XSTEPDOWN_XCORESTATE_XU63 XU63 (
.i0(net_404),
.i1(net_413),
.i2(net_443),
.i3(net_446),
.i4(net_449),
.i5(net_450),
.i6(net_453),
.i7(net_456),
.i8(net_457),
.sr(net_414),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU64 XU64 (
.i0(net_418),
.i1(net_463),
.sr(net_423),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU65 XU65 (
.i0(net_387),
.i1(net_463),
.sr(net_399),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU66 XU66 (
.i0(net_417),
.i1(net_418),
.sr(net_410),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSR2_XU1_XSTEPDOWN_XCORESTATE_XU67 XU67 (
.i0(net_445),
.i1(net_404),
.sr(net_422),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT3_0_XU1_XSTEPDOWN_XCORESTATE_XU68 XU68 (
.o(enable_fault),
.tstate0(net_390),
.tstate1(net_394),
.tstate2(net_405),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT2_0_XU1_XSTEPDOWN_XCORESTATE_XU69 XU69 (
.o(enable_powergood),
.tstate0(net_394),
.tstate1(net_405),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmSTATE8DF_XU1_XSTEPDOWN_XCORESTATE_XU7 XU7 (
.r0(net_389),
.r1(net_414),
.r2(net_423),
.s0(net_399),
.s1(net_410),
.s2(net_422),
.porb(porb),
.state0(net_385),
.state1(net_391),
.state2(net_400),
.state3(net_390),
.state4(net_411),
.state5(net_415),
.state6(net_394),
.state7(net_405),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.hjconfig_0(net_375),
.hjconfig_1(net_376),
.hjconfig_2(net_377),
.hjconfig_3(net_378),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_1_XU1_XSTEPDOWN_XCORESTATE_XU71 XU71 (
.o(enable_softstart),
.i0(ok_regulation),
.tstate(net_405),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XCORESTATE_XU72 XU72 (
.o(enable_discharge),
.tstate(net_391),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT3_0_XU1_XSTEPDOWN_XCORESTATE_XU74 XU74 (
.o(enable_driver),
.tstate0(net_390),
.tstate1(net_394),
.tstate2(net_405),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT1_0_XU1_XSTEPDOWN_XCORESTATE_XU75 XU75 (
.o(fault_core),
.tstate(net_400),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

VESPAasmOUTPUT5_0_XU1_XSTEPDOWN_XCORESTATE_XU9 XU9 (
.o(enable_feedback),
.tstate0(net_390),
.tstate1(net_411),
.tstate2(net_394),
.tstate3(net_405),
.tstate4(net_391),
.CELG59462(CELG59462),
.CELV96848(CELV96848),
.CELSUB40948(CELSUB40948)
);

inv_XU1_XSTEPDOWN_XCORESTATE_XU1 XU1 (
.i(ok_feedback),
.o(net_398),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XCORESTATE_XU2 XU2 (
.i(ok_driver),
.o(net_421),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XCORESTATE_XU3 XU3 (
.i(ok_fault),
.o(net_432),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XCORESTATE_XU4 XU4 (
.i(ok_regulation),
.o(net_439),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XCORESTATE_XU5 XU5 (
.i(ok_powergood),
.o(net_447),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XCORESTATE_XU6 XU6 (
.i(ok_service),
.o(net_436),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU12 XU12 (
.i(net_402),
.o(net_401),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU14 XU14 (
.i(net_424),
.o(net_425),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU15 XU15 (
.i(net_424),
.o(net_429),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU17 XU17 (
.i(net_441),
.o(net_440),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU19 XU19 (
.i(net_455),
.o(net_451),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU20 XU20 (
.i(net_455),
.o(net_454),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU22 XU22 (
.i(net_462),
.o(net_459),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU23 XU23 (
.i(net_462),
.o(net_461),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU25 XU25 (
.i(net_470),
.o(net_466),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU26 XU26 (
.i(net_470),
.o(net_469),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU28 XU28 (
.i(net_477),
.o(net_476),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU30 XU30 (
.i(net_482),
.o(net_479),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

delayfixed_XU1_XSTEPDOWN_XCORESTATE_XU31 XU31 (
.i(net_482),
.o(net_481),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU76 XU76 (
.i(net_385),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_OFF(tdi_STEPDOWNalgorithmCORE0p0_OFF_XU76),
.ten_STEPDOWNalgorithmCORE0p0_OFF(ten_STEPDOWNalgorithmCORE0p0_OFF_XU76)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU77 XU77 (
.i(net_391),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_DISCHARGE(tdi_STEPDOWNalgorithmCORE0p0_DISCHARGE_XU77),
.ten_STEPDOWNalgorithmCORE0p0_DISCHARGE(ten_STEPDOWNalgorithmCORE0p0_DISCHARGE_XU77)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU78 XU78 (
.i(net_400),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_FAULT(tdi_STEPDOWNalgorithmCORE0p0_FAULT_XU78),
.ten_STEPDOWNalgorithmCORE0p0_FAULT(ten_STEPDOWNalgorithmCORE0p0_FAULT_XU78)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU79 XU79 (
.i(net_390),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_POWERUP(tdi_STEPDOWNalgorithmCORE0p0_POWERUP_XU79),
.ten_STEPDOWNalgorithmCORE0p0_POWERUP(ten_STEPDOWNalgorithmCORE0p0_POWERUP_XU79)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU80 XU80 (
.i(net_411),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_POWERDOWN(tdi_STEPDOWNalgorithmCORE0p0_POWERDOWN_XU80),
.ten_STEPDOWNalgorithmCORE0p0_POWERDOWN(ten_STEPDOWNalgorithmCORE0p0_POWERDOWN_XU80)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU81 XU81 (
.i(net_415),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_UNDEF5(tdi_STEPDOWNalgorithmCORE0p0_UNDEF5_XU81),
.ten_STEPDOWNalgorithmCORE0p0_UNDEF5(ten_STEPDOWNalgorithmCORE0p0_UNDEF5_XU81)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU82 XU82 (
.i(net_394),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_RUN(tdi_STEPDOWNalgorithmCORE0p0_RUN_XU82),
.ten_STEPDOWNalgorithmCORE0p0_RUN(ten_STEPDOWNalgorithmCORE0p0_RUN_XU82)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU83 XU83 (
.i(net_405),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_SOFTSTART(tdi_STEPDOWNalgorithmCORE0p0_SOFTSTART_XU83),
.ten_STEPDOWNalgorithmCORE0p0_SOFTSTART(ten_STEPDOWNalgorithmCORE0p0_SOFTSTART_XU83)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU84 XU84 (
.i(enable_fault),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_enable_fault(tdi_STEPDOWNalgorithmCORE0p0_enable_fault_XU84),
.ten_STEPDOWNalgorithmCORE0p0_enable_fault(ten_STEPDOWNalgorithmCORE0p0_enable_fault_XU84)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU85 XU85 (
.i(enable_feedback),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_enable_feedback(tdi_STEPDOWNalgorithmCORE0p0_enable_feedback_XU85),
.ten_STEPDOWNalgorithmCORE0p0_enable_feedback(ten_STEPDOWNalgorithmCORE0p0_enable_feedback_XU85)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU86 XU86 (
.i(enable_powergood),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_enable_powergood(tdi_STEPDOWNalgorithmCORE0p0_enable_powergood_XU86),
.ten_STEPDOWNalgorithmCORE0p0_enable_powergood(ten_STEPDOWNalgorithmCORE0p0_enable_powergood_XU86)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU87 XU87 (
.i(enable_softstart),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_enable_softstart(tdi_STEPDOWNalgorithmCORE0p0_enable_softstart_XU87),
.ten_STEPDOWNalgorithmCORE0p0_enable_softstart(ten_STEPDOWNalgorithmCORE0p0_enable_softstart_XU87)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU88 XU88 (
.i(enable_discharge),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_enable_discharge(tdi_STEPDOWNalgorithmCORE0p0_enable_discharge_XU88),
.ten_STEPDOWNalgorithmCORE0p0_enable_discharge(ten_STEPDOWNalgorithmCORE0p0_enable_discharge_XU88)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU89 XU89 (
.i(enable_regulation),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_enable_regulation(tdi_STEPDOWNalgorithmCORE0p0_enable_regulation_XU89),
.ten_STEPDOWNalgorithmCORE0p0_enable_regulation(ten_STEPDOWNalgorithmCORE0p0_enable_regulation_XU89)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU90 XU90 (
.i(enable_driver),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_enable_driver(tdi_STEPDOWNalgorithmCORE0p0_enable_driver_XU90),
.ten_STEPDOWNalgorithmCORE0p0_enable_driver(ten_STEPDOWNalgorithmCORE0p0_enable_driver_XU90)
);

dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU91 XU91 (
.i(fault_core),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_STEPDOWNalgorithmCORE0p0_fault_core(tdi_STEPDOWNalgorithmCORE0p0_fault_core_XU91),
.ten_STEPDOWNalgorithmCORE0p0_fault_core(ten_STEPDOWNalgorithmCORE0p0_fault_core_XU91)
);

DFTtm8d dft_hex0x5 (
.G(CELG59462),
.V(CELV96848),
.a({a1,a0}),
.SUB(CELSUB40948),
.tdi({tdi_STEPDOWNalgorithmCORE0p0_SOFTSTART_XU83,tdi_STEPDOWNalgorithmCORE0p0_RUN_XU82,tdi_STEPDOWNalgorithmCORE0p0_UNDEF5_XU81,tdi_STEPDOWNalgorithmCORE0p0_POWERDOWN_XU80,tdi_STEPDOWNalgorithmCORE0p0_POWERUP_XU79,tdi_STEPDOWNalgorithmCORE0p0_FAULT_XU78,tdi_STEPDOWNalgorithmCORE0p0_DISCHARGE_XU77,tdi_STEPDOWNalgorithmCORE0p0_OFF_XU76}),
.tdo(tdo),
.ten({ten_STEPDOWNalgorithmCORE0p0_SOFTSTART_XU83,ten_STEPDOWNalgorithmCORE0p0_RUN_XU82,ten_STEPDOWNalgorithmCORE0p0_UNDEF5_XU81,ten_STEPDOWNalgorithmCORE0p0_POWERDOWN_XU80,ten_STEPDOWNalgorithmCORE0p0_POWERUP_XU79,ten_STEPDOWNalgorithmCORE0p0_FAULT_XU78,ten_STEPDOWNalgorithmCORE0p0_DISCHARGE_XU77,ten_STEPDOWNalgorithmCORE0p0_OFF_XU76}),
.tma({a0,a0,a0,a0,a0,a1,a0,a1}),
.tmi(tmi[4:0])
);

DFTtm8d dft_hex0x6 (
.G(CELG59462),
.V(CELV96848),
.a({b1,b0}),
.SUB(CELSUB40948),
.tdi({tdi_STEPDOWNalgorithmCORE0p0_fault_core_XU91,tdi_STEPDOWNalgorithmCORE0p0_enable_driver_XU90,tdi_STEPDOWNalgorithmCORE0p0_enable_regulation_XU89,tdi_STEPDOWNalgorithmCORE0p0_enable_discharge_XU88,tdi_STEPDOWNalgorithmCORE0p0_enable_softstart_XU87,tdi_STEPDOWNalgorithmCORE0p0_enable_powergood_XU86,tdi_STEPDOWNalgorithmCORE0p0_enable_feedback_XU85,tdi_STEPDOWNalgorithmCORE0p0_enable_fault_XU84}),
.tdo(tdo),
.ten({ten_STEPDOWNalgorithmCORE0p0_fault_core_XU91,ten_STEPDOWNalgorithmCORE0p0_enable_driver_XU90,ten_STEPDOWNalgorithmCORE0p0_enable_regulation_XU89,ten_STEPDOWNalgorithmCORE0p0_enable_discharge_XU88,ten_STEPDOWNalgorithmCORE0p0_enable_softstart_XU87,ten_STEPDOWNalgorithmCORE0p0_enable_powergood_XU86,ten_STEPDOWNalgorithmCORE0p0_enable_feedback_XU85,ten_STEPDOWNalgorithmCORE0p0_enable_fault_XU84}),
.tma({b0,b0,b0,b0,b0,b1,b1,b0}),
.tmi(tmi[4:0])
);

drm32 drm_hex0x10 (
.G(CELG59462),
.V(CELV96848),
.d0(d0),
.d1(d1),
.id({d0,d0,d0,d1,d0,d0,d0,d0}),
.SUB(CELSUB40948),
.tmi(tmi[4:0]),
.drm0({net_320,net_319,net_308,net_307,net_306,net_305,net_304,net_303}),
.drm1({net_360,net_359,net_352,net_351,net_336,net_335,net_322,net_321}),
.drm2({net_350,net_349,net_348,net_347,net_346,net_345,net_344,net_343}),
.drm3({noconn_drm32_drm3_7,noconn_drm32_drm3_6,net_378,net_377,net_376,net_375,net_368,net_367}),
.por0({d0,d0,d0,d0,d0,d0,d0,d0}),
.por1({d0,d0,d0,d0,d0,d0,d0,d0}),
.por2({d0,d0,d0,d0,d0,d0,d0,d0}),
.por3({d0,d0,d0,d0,d0,d0,d0,d0}),
.bypload(d0),
.lastdrm(d0)
);

STONEnoconn XNCnoconn_drm32_drm3_6 (
.noconn(noconn_drm32_drm3_6)
);

STONEnoconn XNCnoconn_drm32_drm3_7 (
.noconn(noconn_drm32_drm3_7)
);

endmodule

