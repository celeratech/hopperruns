module dftprobe_XLOOP_XCONTROL_XU72 (i,tdi_STEPDOWNalgorithmCONTROL1p3_botstate,ten_STEPDOWNalgorithmCONTROL1p3_botstate,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_botstate;
input  ten_STEPDOWNalgorithmCONTROL1p3_botstate;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

