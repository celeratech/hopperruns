//Celera:levelshifter0L2H_fetdriver_XLOOP_XDRIVER_XTOPDRIVER_XTSWDRIVER_Xfetin
//Celera Confidential Symbol Generator
//Direction: low2high, Maximum high voltage:36V 
//Enable pin:yes
module levelshifter0L2H_fetdriver_XLOOP_XDRIVER_XTOPDRIVER_XTSWDRIVER_Xfetin (SIMPV,CELSUB,HVPOS,HVNEG,in,out,
enable_levelshifter,
CELG);
input SIMPV;
input CELG;
input CELSUB;
input HVPOS;
input HVNEG;
input in;
output out;
input enable_levelshifter;
endmodule

