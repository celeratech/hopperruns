module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU41 (i,tdi_SOFTSTARTinternalNOFAULT_enable_startup,ten_SOFTSTARTinternalNOFAULT_enable_startup,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTinternalNOFAULT_enable_startup;
input  ten_SOFTSTARTinternalNOFAULT_enable_startup;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

