//Celera:voltage2current_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU3
//Celera Confidential Symbol Generator
//Gain: 25, Direction: source, Iout Clamp: no
//DFT:no, Accuracy: na, Input Stage Type: na
module voltage2current_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU3 (CELV,SUB,enable_voltage2current,IP,ok_voltage2current,IOUT,VIN,ten,
CELG);
input CELV;
input SUB;
input enable_voltage2current;
input IP;
output ok_voltage2current;
output IOUT;
input VIN;
input ten;
input CELG;
endmodule

