//Celera:delay0_delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU3_XU20_delay0
//TYPE:fixed 5us EDGE:rise DFT:no ACC:no
module delay0_delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU3_XU20_delay0 (i,CELV,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELSUB;
input CELG;
endmodule

