//Celera:inv_XU1_XSERVICE_XU14_XU3
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSERVICE_XU14_XU3 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

