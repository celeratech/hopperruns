module dfthijack_XU1_XSTEPDOWN_XDISCHARGE_XU4_XU4 (HIJACKdischargeo,CELG,CELV,CELSUB,ten_HIJACKdischargeenable,ten_HIJACKdischargestatus,HIJACKdischarge);
output  HIJACKdischargeo;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HIJACKdischargeenable;
input  ten_HIJACKdischargestatus;
input  HIJACKdischarge;
endmodule

