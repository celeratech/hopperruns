//Celera:porb_XU1_XSERVICE_XBIASSERVICE_XU9
//Global PORB
module porb_XU1_XSERVICE_XBIASSERVICE_XU9 (CELV,SENSE_PORB,porb,
enable_porb,CELG,SUB);
input CELV;
input SENSE_PORB;
output porb;
input enable_porb;
input SUB;
input CELG;
endmodule

