module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU36 (i,tdi_SOFTSTARTinternalNOFAULT_STARTUP,ten_SOFTSTARTinternalNOFAULT_STARTUP,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTinternalNOFAULT_STARTUP;
input  ten_SOFTSTARTinternalNOFAULT_STARTUP;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

