module dftprobe_XU1_XSTEPDOWN_XFAULT_XU1_XU9 (i,tdi_FAULTdetect,ten_FAULTdetect,CELG,CELSUB,CELV);
input  i;
output  tdi_FAULTdetect;
input  ten_FAULTdetect;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

