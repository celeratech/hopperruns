//Celera:nor3_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU9_XU11
//Celera Confidential Symbol Generator
//NOR3
module nor3_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU9_XU11 (CELV,CELG,i0,i1,i2,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input i2;
input SUB;
output o;
endmodule

