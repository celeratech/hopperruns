//Celera:oneshot_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU2
//Celera Confidential Symbol Generator
//One Shot50ns OneShot - Bad Designer!!
module oneshot_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU2 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

