//Celera:timingskew_XLOOP_XCONTROL_XU38_XU10
//Celera Confidential Symbol Generator
//TYPE:rise Bits:2 with 2.0ns LSB
module timingskew_XLOOP_XCONTROL_XU38_XU10 (CELV,in,out,
s,
CELG,CELSUB);
input CELV;
input in;
output out;
input [1:0] s;
input CELG;
input CELSUB;
endmodule

