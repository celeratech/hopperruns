//Celera:dbuf_XLOOP_XDRIVER_XTOPDRIVER_XU23
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XLOOP_XDRIVER_XTOPDRIVER_XU23 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

