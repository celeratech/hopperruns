module dfthijack_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU4 (HJregulationeno,CELG,CELV,CELSUB,ten_HJregulationenenable,ten_HJregulationenstatus,HJregulationen);
output  HJregulationeno;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJregulationenenable;
input  ten_HJregulationenstatus;
input  HJregulationen;
endmodule

