module dftprobe_XLOOP_XREG_XDEBUG_XU13 (i,TAI_REGiref,ten_REGiref,CELG,CELSUB,CELV);
input  i;
output  TAI_REGiref;
input  ten_REGiref;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

