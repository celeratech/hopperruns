//Celera:logicshifter0L2H_fetdriver_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWDRIVE_Xglobal
//Logic Level shifter with Enable
module logicshifter0L2H_fetdriver_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWDRIVE_Xglobal (enable_logicshifter,
VIN1,VIN2,
in,
out,
CELG,CELSUB);
input VIN1;
input VIN2;
input in;
output out;
input enable_logicshifter;
input CELSUB;
input CELG;
endmodule

