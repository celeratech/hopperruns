//Celera:capacitorfixed_XLOOP_XREG_XFREQ_XU27
//Celera Confidential Symbol Generator
//CAPACITOR CONTROL:capacitor
//VALUE: 30.00pF TYPE:mim
module capacitorfixed_XLOOP_XREG_XFREQ_XU27 (CP,
CN);
inout CP;
inout CN;
endmodule

