//Celera:capacitorfixed_slopecomp_XLOOP_XDRIVER_XTOPSW_XU38_Xslc
//Celera Confidential Symbol Generator
//CAPACITOR CONTROL:capacitor
//VALUE: 15.00pF TYPE:mim
module capacitorfixed_slopecomp_XLOOP_XDRIVER_XTOPSW_XU38_Xslc (CP,
CN);
inout CP;
inout CN;
endmodule

