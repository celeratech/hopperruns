//Celera:levelshifter0H2L_XLOOP_XDRIVER_XTOPDRIVER_XU7
//Celera Confidential Symbol Generator
//Direction: high2low, Maximum high voltage:36V 
//Enable pin:no
module levelshifter0H2L_XLOOP_XDRIVER_XTOPDRIVER_XU7 (SIMPV,CELSUB,HVPOS,HVNEG,in,out,
CELG);
input SIMPV;
input CELG;
input CELSUB;
input HVPOS;
input HVNEG;
input in;
output out;
endmodule

