module dftprobe_XU1_XSERVICE_XATESERVICE_XU21 (i,tdi_encore,ten_encore,CELG,CELSUB,CELV);
input  i;
output  tdi_encore;
input  ten_encore;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

