module dftprobe_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU1 (i,tdi_POWERGOODstartup,ten_POWERGOODstartup,CELG,CELSUB,CELV);
input  i;
output  tdi_POWERGOODstartup;
input  ten_POWERGOODstartup;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

