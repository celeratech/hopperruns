//Celera:delayfixed_XLOOP_XCONTROL_XU11_XU6
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:rise
module delayfixed_XLOOP_XCONTROL_XU11_XU6 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

