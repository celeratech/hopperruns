//Celera:nor4_XLOOP_XCONTROL_XU34_XU18
//Celera Confidential Symbol Generator
//nor4
module nor4_XLOOP_XCONTROL_XU34_XU18 (CELV,CELG,i0,i1,i2,i3,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input i2;
input i3;
input SUB;
output o;
endmodule

