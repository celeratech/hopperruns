module dfthijack_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU10 (POWGOODoutputo,CELG,CELV,CELSUB,ten_POWGOODoutputenable,ten_POWGOODoutputstatus,POWGOODoutput);
output  POWGOODoutputo;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_POWGOODoutputenable;
input  ten_POWGOODoutputstatus;
input  POWGOODoutput;
endmodule

