module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU88 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_discharge,ten_STEPDOWNalgorithmCORE0p0_enable_discharge,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_enable_discharge;
input  ten_STEPDOWNalgorithmCORE0p0_enable_discharge;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

