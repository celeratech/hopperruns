module dftprobe_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU18 (i,tdi_botswzcross,ten_botswzcross,CELG,CELSUB,CELV);
input  i;
output  tdi_botswzcross;
input  ten_botswzcross;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

