module dfthijack_XU1_XSTEPDOWN_XSOFTSTART_XU7_XU9 (ENABLEsoftstarto,CELG,CELV,CELSUB,ten_ENABLEsoftstartenable,ten_ENABLEsoftstartstatus,ENABLEsoftstart);
output  ENABLEsoftstarto;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_ENABLEsoftstartenable;
input  ten_ENABLEsoftstartstatus;
input  ENABLEsoftstart;
endmodule

