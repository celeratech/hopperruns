module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU75 (i,tdi_STEPDOWNalgorithmCONTROL0p2_IDLE,ten_STEPDOWNalgorithmCONTROL0p2_IDLE,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_IDLE;
input  ten_STEPDOWNalgorithmCONTROL0p2_IDLE;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

