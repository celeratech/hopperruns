module dfthijack_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU20 (hjenable_drivero,CELG,CELV,CELSUB,ten_hjenable_driverenable,ten_hjenable_driverstatus,hjenable_driver);
output  hjenable_drivero;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_hjenable_driverenable;
input  ten_hjenable_driverstatus;
input  hjenable_driver;
endmodule

