//Celera:dbuf_XU1_XSTEPDOWN_XCORESTATE_XU75_XU25
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XCORESTATE_XU75_XU25 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

