//Celera:tie_XU1_XSERVICE_XATESERVICE_XU15
//Celera Confidential Symbol Generator
//TIE
module tie_XU1_XSERVICE_XATESERVICE_XU15 (CELV,CELG,a1,SUB);
input CELV;
input CELG;
output a1;
input SUB;
endmodule

