module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU90 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_driver,ten_STEPDOWNalgorithmCORE0p0_enable_driver,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_enable_driver;
input  ten_STEPDOWNalgorithmCORE0p0_enable_driver;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

