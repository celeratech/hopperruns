//Celera:dbuf_XU1_XSTEPDOWN_XSOFTSTART_XU8_XU16_XU19
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XSOFTSTART_XU8_XU16_XU19 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

