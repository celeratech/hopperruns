module dftprobe_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU17 (i,TAI_REGULATIONiref,ten_REGULATIONiref,CELG,CELSUB,CELV);
input  i;
output  TAI_REGULATIONiref;
input  ten_REGULATIONiref;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

