//Celera:fet_fet_XLOOP_XDRIVER_XTOPDRIVER_XTOPSW_Xfet
//Celera Confidential Symbol Generator
//power NMOS:Ron:0.100 Ohm
//Vgs 6V Vds 6V
//Kelvin:no

module fet_fet_XLOOP_XDRIVER_XTOPDRIVER_XTOPSW_Xfet (GATE,SOURCE,DRAIN,NMOSiso6,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
input NMOSiso6;
endmodule

