//Celera:fet_fetdriver_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWDRIVE_Xpmos0
//Celera Confidential Symbol Generator
//power PMOS:Ron:2.000 Ohm
//Vgs 6V Vds 6V
//Kelvin:no

module fet_fetdriver_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWDRIVE_Xpmos0 (GATE,DRAIN,
SOURCE,
PMOSiso6,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
input PMOSiso6;
endmodule

