module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU83 (i,tdi_STEPDOWNalgorithmCORE0p0_SOFTSTART,ten_STEPDOWNalgorithmCORE0p0_SOFTSTART,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_SOFTSTART;
input  ten_STEPDOWNalgorithmCORE0p0_SOFTSTART;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

