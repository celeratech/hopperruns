//Celera:dbuf_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU7
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XPOWERGOOD_XU6_XU7 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

