//Celera:celeradacr2r_XU1_XSTEPDOWN_XSOFTSTART_XU9_XU5
//Celera Confidential Symbol Generator
//LADDER DAC:6 Bits 500.0K with output Buffer
module celeradacr2r_XU1_XSTEPDOWN_XSOFTSTART_XU9_XU5 (SIMPV,
global_dac,DAC,ok_dac,
IP,
i,
strobe_dac,
DACREF,
GNDSENSE,
CELG,CELSUB); 
input SIMPV;
input DACREF;
input global_dac;
output DAC;
input strobe_dac;
output ok_dac;
input IP;
input [5:0] i;
input GNDSENSE;
input CELG;
input CELSUB;
endmodule

