//Celera:delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU31_XU3
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:both
module delayfixed_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU31_XU3 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

