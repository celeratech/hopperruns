//Celera:fet_fet_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xnmos0_Xfet
//Celera Confidential Symbol Generator
//power NMOS:Ron:2.000 Ohm
//Vgs 6V Vds 6V
//Kelvin:no

module fet_fet_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xnmos0_Xfet (GATE,SOURCE,DRAIN,NMOSiso6,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
input NMOSiso6;
endmodule

