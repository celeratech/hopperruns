//Celera:resistordivider_XLOOP_XREGULATION_XU2_XU23
//Celera Confidential Symbol Generator
//VMAX:6V R:1000.0KOhm 1Taps
module resistordivider_XLOOP_XREGULATION_XU2_XU23 (TOP,
TAP0,
CELG, BOTTOM);
inout TOP;
output TAP0;
input CELG;
inout BOTTOM;
endmodule

