module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU7_XU2 (i,tdi_SOFTSTARTtime,ten_SOFTSTARTtime,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTtime;
input  ten_SOFTSTARTtime;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

