module dftprobe_XU1_XSERVICE_XATESERVICE_XU4 (i,tdi_ok_mudv,ten_ok_mudv,CELG,CELSUB,CELV);
input  i;
output  tdi_ok_mudv;
input  ten_ok_mudv;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

