module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU42 (i,tdi_SOFTSTARTinternalNOFAULT_enable_charge,ten_SOFTSTARTinternalNOFAULT_enable_charge,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTinternalNOFAULT_enable_charge;
input  ten_SOFTSTARTinternalNOFAULT_enable_charge;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

