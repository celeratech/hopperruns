//Celera:dbuf_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU28
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU28 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

