//Celera:nor3_XLOOP_XCONTROL_XU55_XU2
//Celera Confidential Symbol Generator
//NOR3
module nor3_XLOOP_XCONTROL_XU55_XU2 (CELV,CELG,i0,i1,i2,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input i2;
input SUB;
output o;
endmodule

