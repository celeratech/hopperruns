module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU86 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_powergood,ten_STEPDOWNalgorithmCORE0p0_enable_powergood,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_enable_powergood;
input  ten_STEPDOWNalgorithmCORE0p0_enable_powergood;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

