module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU40 (i,tdi_SOFTSTARTinternalNOFAULT_state_off,ten_SOFTSTARTinternalNOFAULT_state_off,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTinternalNOFAULT_state_off;
input  ten_SOFTSTARTinternalNOFAULT_state_off;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

