module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU69 (i,tdi_STEPDOWNalgorithmCONTROL0p2_OFF,ten_STEPDOWNalgorithmCONTROL0p2_OFF,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_OFF;
input  ten_STEPDOWNalgorithmCONTROL0p2_OFF;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

