//Celera:timingskew_XLOOP_XDRIVER_XBBMDRIVER_XU14
//Celera Confidential Symbol Generator
//TYPE:fall Bits:5 with 2.0ns LSB
module timingskew_XLOOP_XDRIVER_XBBMDRIVER_XU14 (CELV,in,out,
factory_timingskew,
CELG,CELSUB);
input CELV;
input in;
output out;
input [4:0] factory_timingskew;
input CELG;
input CELSUB;
endmodule

