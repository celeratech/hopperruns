//Celera:padopendrain_XU1_XSTEPDOWN_XPOWERGOOD_XU10_XU2
//Celera Confidential Symbol Generator
//Open Drain output PAD with 6V, Ron 50 Ohms
//No Glitch filter
//ON Logic:invert polarity
//DFT:no TESTMODE:no RETURN PIN:no
module padopendrain_XU1_XSTEPDOWN_XPOWERGOOD_XU10_XU2 (CELV, input_padopendrain, PAD, 
CELG, SUB ); 
input CELV;
input input_padopendrain;
input CELG;
input SUB;
inout PAD;
endmodule

