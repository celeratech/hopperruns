module dftprobe_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU38 (i,tdi_SOFTSTARTinternalNOFAULT_CHARGE,ten_SOFTSTARTinternalNOFAULT_CHARGE,CELG,CELSUB,CELV);
input  i;
output  tdi_SOFTSTARTinternalNOFAULT_CHARGE;
input  ten_SOFTSTARTinternalNOFAULT_CHARGE;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

