//Celera:inv_XU1_XSERVICE_XBIASSERVICE_XU8
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSERVICE_XBIASSERVICE_XU8 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

