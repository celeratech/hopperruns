module dfthijack_XLOOP_XDRIVER_XDEBUG_XU6 (HJdrvbso,CELG,CELV,CELSUB,ten_HJdrvbsenable,ten_HJdrvbsstatus,HJdrvbs);
output  HJdrvbso;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJdrvbsenable;
input  ten_HJdrvbsstatus;
input  HJdrvbs;
endmodule

