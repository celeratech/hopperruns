//Celera:nor2_XLOOP_XDRIVER_XBBM_XU20
//Celera Confidential Symbol Generator
//nor2
module nor2_XLOOP_XDRIVER_XBBM_XU20 (CELV,CELG,i0,i1,o,SUB);
input CELV;
input CELG;
input i0;
input i1;
input SUB;
output o;
endmodule

