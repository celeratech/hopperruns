//Celera:logicshifter0L2H_fetdriver_XLOOP_XDRIVER_XTOPDRIVER_XTSWDRIVER_Xenable
//Logic Level shifter with Enable
module logicshifter0L2H_fetdriver_XLOOP_XDRIVER_XTOPDRIVER_XTSWDRIVER_Xenable (enable_logicshifter,
HVPOS,HVNEG,SIMPV,
in,
out,
CELG,CELSUB);
input HVPOS;
input HVNEG;
input SIMPV;
input in;
output out;
input enable_logicshifter;
input CELSUB;
input CELG;
endmodule

