module dftprobe_XLOOP_XDRIVER_XDEBUG_XU11 (i,tdi_DRVtopswstatus,ten_DRVtopswstatus,CELG,CELSUB,CELV);
input  i;
output  tdi_DRVtopswstatus;
input  ten_DRVtopswstatus;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

