module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU76 (i,tdi_STEPDOWNalgorithmCORE0p0_OFF,ten_STEPDOWNalgorithmCORE0p0_OFF,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_OFF;
input  ten_STEPDOWNalgorithmCORE0p0_OFF;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

