//Celera:resistordivider_vbias_XU1_XSERVICE_XBIASSERVICE_XU1_XRuvlo
//Celera Confidential Symbol Generator
//VMAX:6V R:6000.0KOhm 1Taps
module resistordivider_vbias_XU1_XSERVICE_XBIASSERVICE_XU1_XRuvlo (TOP,
TAP0,
CELG, BOTTOM);
inout TOP;
output TAP0;
input CELG;
inout BOTTOM;
endmodule

