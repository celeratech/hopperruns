module dfthijack_XU1_XSTEPDOWN_XFAULT_XU1_XU6 (HIJACKfaultENABLEo,CELG,CELV,CELSUB,ten_HIJACKfaultENABLEenable,ten_HIJACKfaultENABLEstatus,HIJACKfaultENABLE);
output  HIJACKfaultENABLEo;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HIJACKfaultENABLEenable;
input  ten_HIJACKfaultENABLEstatus;
input  HIJACKfaultENABLE;
endmodule

