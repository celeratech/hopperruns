//Celera:bgcomp_XU1_XSERVICE_XBIASSERVICE_XU4
//Celera Confidential Symbol Generator
//Trip threshold: 1.2V, Maximum Supply Voltage: 30V, Maximum Input Voltage:30V
//Logic shift output:yes, Trim trip threshold: yes, Enable pin: no, DFT: no
module bgcomp_XU1_XSERVICE_XBIASSERVICE_XU4 (CELSUB,CELPOS,IN,out,global_bgcomp,
CELV,
trim_bgcomp,
CELG);
input CELSUB;
input CELPOS;
input IN;
output out;
input global_bgcomp;
input CELV;
input [7:0] trim_bgcomp;
input CELG;
endmodule

