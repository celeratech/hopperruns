//Celera:inv_XU1_XSTEPDOWN_XCORESTATE_XU21_XU9
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSTEPDOWN_XCORESTATE_XU21_XU9 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

