// ------------------------ Module Definitions -----------
module dbufdft_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14 (i,o,CELG,CELV,CELSUB,tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14,ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf0,ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf1);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14;
  input  ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf0;
  input  ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf1;
endmodule

module dbufdft_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28 (i,o,CELG,CELV,CELSUB,tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28,ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf0,ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf1);
  input  i;
  output  o;
  input  CELG;
  input  CELV;
  input  CELSUB;
  output  tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28;
  input  ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf0;
  input  ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf1;
endmodule

module nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU2 (CELV,CELG,i0,i1,i2,o,SUB);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module dff_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU8 (CELV,CELG,d,rb,ck,q,qb,SUB);
  input  d;
  output  q;
  input  ck;
  output  qb;
  input  rb;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module tie_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU9 (CELV,CELG,a1,SUB);
  output  a1;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU11 (CELV,in,out,factory_timingskew,CELG,CELSUB);
  input  in;
  output  out;
  input  CELG;
  input  CELV;
  input  CELSUB;
  input [4:0] factory_timingskew;
endmodule

module nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU12 (CELV,CELG,i0,i1,i2,o,SUB);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU15 (CELV,in,out,factory_timingskew,CELG,CELSUB);
  input  in;
  output  out;
  input  CELG;
  input  CELV;
  input  CELSUB;
  input [4:0] factory_timingskew;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU16 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU17 (CELV,CELG,i0,i1,i2,o,SUB);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU18 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU19 (CELV,CELG,i0,i1,i2,o,SUB);
  output  o;
  input  i0;
  input  i1;
  input  i2;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU20 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU21 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module nor2_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU22 (CELV,CELG,i0,i1,o,SUB);
  output  o;
  input  i0;
  input  i1;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU24 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU25 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module nor2_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU26 (CELV,CELG,i0,i1,o,SUB);
  output  o;
  input  i0;
  input  i1;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module dff_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU27 (CELV,CELG,d,rb,ck,q,qb,SUB);
  input  d;
  output  q;
  input  ck;
  output  qb;
  input  rb;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU30 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU33 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU38 (CELV,in,out,factory_timingskew,CELG,CELSUB);
  input  in;
  output  out;
  input  CELG;
  input  CELV;
  input  CELSUB;
  input [4:0] factory_timingskew;
endmodule

module tie_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU39 (CELV,CELG,a1,SUB);
  output  a1;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

module timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU41 (CELV,in,out,factory_timingskew,CELG,CELSUB);
  input  in;
  output  out;
  input  CELG;
  input  CELV;
  input  CELSUB;
  input [4:0] factory_timingskew;
endmodule

module inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU47 (CELV,CELG,i,o,SUB);
  input  i;
  output  o;
  input  SUB;
  input  CELG;
  input  CELV;
endmodule

//Verilog HDL for "Generate", "STONEnoconn" "functional"


module STONEnoconn ( noconn );

  input noconn;
endmodule


module fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWIREP (GATE,SOURCE,DRAIN,SOURCEk,DRAINk,IREPLICA,SUB);
  input  SUB;
  input  GATE;
  inout  DRAIN;
  inout  DRAINk;
  inout  SOURCE;
  inout  SOURCEk;
  inout  IREPLICA;
endmodule

module currentlimitfet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZERO (SIMPV,SUB,measure_currentlimit,VSENSE,IREPLICA,currentlimit,enable_currentlimit,trim_currentlimit,factory_currentlimit_blanking,IP,global_currentlimit,ten_currentlimit,ten_taext_currentlimit,ten_measure_currentlimit,TAEXT_CURRENTLIMIT,tdi_currentlimit,tdi_currentlimitlive,ten_currentlimit_delay,CELG);
  input  IP;
  input  SUB;
  input  CELG;
  input  SIMPV;
  input  VSENSE;
  input  IREPLICA;
  output  currentlimit;
  output  tdi_currentlimit;
  input  ten_currentlimit;
  input [7:0] trim_currentlimit;
  input  TAEXT_CURRENTLIMIT;
  input  enable_currentlimit;
  input  global_currentlimit;
  input  measure_currentlimit;
  output  tdi_currentlimitlive;
  input [4:0] ten_currentlimit_delay;
  input  ten_taext_currentlimit;
  input  ten_measure_currentlimit;
  input [4:0] factory_currentlimit_blanking;
endmodule

module fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZREP (GATE,SOURCE,DRAIN,SOURCEk,DRAINk,IREPLICA,SUB);
  input  SUB;
  input  GATE;
  inout  DRAIN;
  inout  DRAINk;
  inout  SOURCE;
  inout  SOURCEk;
  inout  IREPLICA;
endmodule

//Verilog HDL for "DFT", "DFTtm8d" "functional"


module DFTtm8d ( a, ten, tdo, tmi, G, SUB, V, tdi, tma );

  input V;
  input  [7:0] tma;
  output  [7:0] ten;
  output  [1:0] a;
  inout tdo;
  input  [7:0] tdi;
  input G;
  input SUB;
  inout  [4:0] tmi;
endmodule


//Verilog HDL for "DFT", "DFTtm8t" "functional"


module DFTtm8t ( a, ten, tmi, G, SUB, V, tma );

  input V;
  input  [7:0] tma;
  output  [7:0] ten;
  output  [1:0] a;
  input G;
  input SUB;
  inout  [4:0] tmi;
endmodule


//Verilog HDL for "DRM", "drm56" "functional"


module drm56 ( V, G, SUB, tmi, bypload, lastdrm, id, por0, por1, por2, por3,
por4, por5, por6, drm0, drm1, drm2, drm3, drm4, drm5, drm6, d1, d0 );

  output  [7:0] drm4;
  input  [7:0] por6;
  input lastdrm;
  input V;
  output d1;
  input  [7:0] por3;
  output  [7:0] drm3;
  input  [7:0] por5;
  input  [7:0] id;
  output d0;
  output  [7:0] drm5;
  output  [7:0] drm2;
  input  [7:0] por2;
  input  [7:0] por1;
  input  [7:0] por4;
  input bypload;
  output  [7:0] drm6;
  output  [7:0] drm0;
  input  [7:0] por0;
  input G;
  output  [7:0] drm1;
  inout  [4:0] tmi;
  input SUB;
endmodule


//Verilog HDL for "DRM", "drm16L" "functional"


module drm16L ( V, G, SUB, tmi, bypload, lastdrm, id, drm0, drm1, d1, d0 );

  input lastdrm;
  input V;
  output d1;
  input  [7:0] id;
  output d0;
  input bypload;
  output  [7:0] drm0;
  input G;
  output  [7:0] drm1;
  inout  [4:0] tmi;
  input SUB;
endmodule


module fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWDRIVER (HVPOS,enable_fetdriverhv,global_fetdriver,fetin,GATE,gate_status,factory_fetdriver_statusadjust,CELG,SIMPV,HVNEG,CELSUB);
  input  CELG;
  output  GATE;
  input  HVNEG;
  input  HVPOS;
  input  SIMPV;
  input  fetin;
  input  CELSUB;
  output  gate_status;
  input  global_fetdriver;
  input  enable_fetdriverhv;
  input [4:0] factory_fetdriver_statusadjust;
endmodule

module currentlimitfet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWCURRENT (SIMPV,SUB,measure_currentlimit,VSENSE,IREPLICA,currentlimit,enable_currentlimit,trim_currentlimit,factory_currentlimit_blanking,IP,global_currentlimit,ten_currentlimit,ten_taext_currentlimit,ten_measure_currentlimit,TAEXT_CURRENTLIMIT,tdi_currentlimit,tdi_currentlimitlive,ten_currentlimit_delay,CELG);
  input  IP;
  input  SUB;
  input  CELG;
  input  SIMPV;
  input  VSENSE;
  input  IREPLICA;
  output  currentlimit;
  output  tdi_currentlimit;
  input  ten_currentlimit;
  input [7:0] trim_currentlimit;
  input  TAEXT_CURRENTLIMIT;
  input  enable_currentlimit;
  input  global_currentlimit;
  input  measure_currentlimit;
  output  tdi_currentlimitlive;
  input [4:0] ten_currentlimit_delay;
  input  ten_taext_currentlimit;
  input  ten_measure_currentlimit;
  input [4:0] factory_currentlimit_blanking;
endmodule

// ------------------------ Module Verilog ---------------
module MUDbotswnmosSdIlimAugment_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2 (SW, tdo, tmi, MUDV, PMUDG, PMUDV, TAEXT, botswon, CELG59462, CELV96848, botswipeak, CELSUB40948, botswstatus, botswzcross, enable_driver, IP_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZERO, IP_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWCURRENT);
inout  SW;
inout  tdo;
inout [4:0] tmi;
input  MUDV;
inout  PMUDG;
input  PMUDV;
input  TAEXT;
input  botswon;
input  CELG59462;
input  CELV96848;
output  botswipeak;
input  CELSUB40948;
output  botswstatus;
output  botswzcross;
input  enable_driver;
input  IP_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZERO;
input  IP_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWCURRENT;


// ------------------------ Wires ------------------------
wire [4:0] tmi;
wire [4:0] factory_timingskew;
wire [7:0] trim_currentlimit;
wire [4:0] ten_currentlimit_delay;
wire [4:0] factory_currentlimit_blanking;
wire [1:0] a;
wire [7:0] tdi;
wire [7:0] ten;
wire [7:0] tma;
wire [7:0] id;
wire [7:0] drm0;
wire [7:0] drm1;
wire [7:0] drm2;
wire [7:0] drm3;
wire [7:0] drm4;
wire [7:0] drm5;
wire [7:0] drm6;
wire [7:0] por0;
wire [7:0] por1;
wire [7:0] por2;
wire [7:0] por3;
wire [7:0] por4;
wire [7:0] por5;
wire [7:0] por6;
wire [4:0] factory_fetdriver_statusadjust;

// ------------------------ Networks ---------------------
dbufdft_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14 XU14 (
.i(net_40),
.o(botswzcross),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14(tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_XU14),
.ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf0(ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf0_XU14),
.ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf1(ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf1_XU14)
);

dbufdft_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28 XU28 (
.i(net_66),
.o(botswipeak),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28(tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_XU28),
.ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf0(ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf0_XU28),
.ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf1(ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf1_XU28)
);

nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU2 XU2 (
.o(net_68),
.i0(net_64),
.i1(net_70),
.i2(net_60),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

dff_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU8 XU8 (
.d(net_45),
.q(net_46),
.ck(net_34),
.qb(net_49),
.rb(net_57),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

tie_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU9 XU9 (
.a1(net_45),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU11 XU11 (
.in(botswstatus),
.out(net_33),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.factory_timingskew({XU11_factory_timingskew_4,XU11_factory_timingskew_3,XU11_factory_timingskew_2,XU11_factory_timingskew_1,XU11_factory_timingskew_0})
);

nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU12 XU12 (
.o(net_61),
.i0(net_59),
.i1(net_63),
.i2(net_60),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU15 XU15 (
.in(botswstatus),
.out(net_59),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.factory_timingskew({XU15_factory_timingskew_4,XU15_factory_timingskew_3,XU15_factory_timingskew_2,XU15_factory_timingskew_1,XU15_factory_timingskew_0})
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU16 XU16 (
.i(net_42),
.o(net_41),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU17 XU17 (
.o(net_42),
.i0(net_38),
.i1(net_46),
.i2(net_34),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU18 XU18 (
.i(net_37),
.o(net_38),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

nand3_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU19 XU19 (
.o(net_35),
.i0(net_33),
.i1(net_37),
.i2(net_34),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU20 XU20 (
.i(net_35),
.o(net_36),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU21 XU21 (
.i(net_39),
.o(net_40),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

nor2_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU22 XU22 (
.o(net_39),
.i0(net_36),
.i1(net_41),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU24 XU24 (
.i(net_68),
.o(net_67),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU25 XU25 (
.i(net_63),
.o(net_64),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

nor2_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU26 XU26 (
.o(net_65),
.i0(net_62),
.i1(net_67),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

dff_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU27 XU27 (
.d(net_69),
.q(net_70),
.ck(net_60),
.qb(net_72),
.rb(net_77),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU30 XU30 (
.i(net_65),
.o(net_66),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU33 XU33 (
.i(net_61),
.o(net_62),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU38 XU38 (
.in(net_33),
.out(net_57),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.factory_timingskew({XU38_factory_timingskew_4,XU38_factory_timingskew_3,XU38_factory_timingskew_2,XU38_factory_timingskew_1,XU38_factory_timingskew_0})
);

tie_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU39 XU39 (
.a1(net_69),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

timingskew_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU41 XU41 (
.in(net_59),
.out(net_77),
.CELG(CELG59462),
.CELV(CELV96848),
.CELSUB(CELSUB40948),
.factory_timingskew({XU41_factory_timingskew_4,XU41_factory_timingskew_3,XU41_factory_timingskew_2,XU41_factory_timingskew_1,XU41_factory_timingskew_0})
);

inv_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU47 XU47 (
.i(net_48),
.o(net_34),
.SUB(CELSUB40948),
.CELG(CELG59462),
.CELV(CELV96848)
);

STONEnoconn XNC43 (
.noconn(net_43)
);

STONEnoconn XNC44 (
.noconn(net_44)
);

STONEnoconn XNC49 (
.noconn(net_49)
);

STONEnoconn XNC72 (
.noconn(net_72)
);

fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWIREP XBOTSWIREP (
.SUB(CELSUB40948),
.GATE(net_56),
.DRAIN(SW),
.DRAINk(net_44),
.SOURCE(PMUDG),
.SOURCEk(net_112),
.IREPLICA(net_111)
);

currentlimitfet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZERO XBOTSWZERO (
.IP(IP_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZERO),
.SUB(CELSUB40948),
.CELG(CELG59462),
.SIMPV(MUDV),
.VSENSE(net_107),
.IREPLICA(net_109),
.currentlimit(net_48),
.tdi_currentlimit(tdi_currentlimit_XBOTSWZERO),
.ten_currentlimit(ten_currentlimit_XBOTSWZERO),
.trim_currentlimit({XBOTSWZERO_trim_currentlimit_7,XBOTSWZERO_trim_currentlimit_6,XBOTSWZERO_trim_currentlimit_5,XBOTSWZERO_trim_currentlimit_4,XBOTSWZERO_trim_currentlimit_3,XBOTSWZERO_trim_currentlimit_2,XBOTSWZERO_trim_currentlimit_1,XBOTSWZERO_trim_currentlimit_0}),
.TAEXT_CURRENTLIMIT(TAEXT),
.enable_currentlimit(enable_driver),
.global_currentlimit(global_currentlimit_XBOTSWZERO),
.measure_currentlimit(botswstatus),
.tdi_currentlimitlive(tdi_currentlimitlive_XBOTSWZERO),
.ten_currentlimit_delay({ten_currentlimit_delay_XBOTSWZERO_4,ten_currentlimit_delay_XBOTSWZERO_3,ten_currentlimit_delay_XBOTSWZERO_2,ten_currentlimit_delay_XBOTSWZERO_1,ten_currentlimit_delay_XBOTSWZERO_0}),
.ten_taext_currentlimit(ten_taext_currentlimit_XBOTSWZERO),
.ten_measure_currentlimit(ten_measure_currentlimit_XBOTSWZERO),
.factory_currentlimit_blanking({XBOTSWZERO_factory_currentlimit_blanking_4,XBOTSWZERO_factory_currentlimit_blanking_3,XBOTSWZERO_factory_currentlimit_blanking_2,XBOTSWZERO_factory_currentlimit_blanking_1,XBOTSWZERO_factory_currentlimit_blanking_0})
);

fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZREP XBOTSWZREP (
.SUB(CELSUB40948),
.GATE(net_56),
.DRAIN(SW),
.DRAINk(net_43),
.SOURCE(PMUDG),
.SOURCEk(net_107),
.IREPLICA(net_109)
);

DFTtm8d dft_hex0x14 (
.G(CELG59462),
.V(CELV96848),
.a({a1,a0}),
.SUB(CELSUB40948),
.tdi({a0,a0,tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_XU28,tdi_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_XU14,tdi_currentlimitlive_XBOTSWZERO,tdi_currentlimit_XBOTSWZERO,tdi_currentlimitlive_XBOTSWCURRENT,tdi_currentlimit_XBOTSWCURRENT}),
.tdo(tdo),
.ten({ten_taext_currentlimit_XBOTSWCURRENT,ten_currentlimit_delay_XBOTSWCURRENT_0,ten_currentlimit_delay_XBOTSWCURRENT_1,ten_currentlimit_delay_XBOTSWCURRENT_2,ten_currentlimit_delay_XBOTSWCURRENT_3,ten_currentlimit_delay_XBOTSWCURRENT_4,global_currentlimit_XBOTSWCURRENT,ten_currentlimit_XBOTSWCURRENT}),
.tma({a0,a0,a0,a1,a0,a1,a0,a0}),
.tmi(tmi[4:0])
);

DFTtm8t dft_hex0x15 (
.G(CELG59462),
.V(CELV96848),
.a({b1,b0}),
.SUB(CELSUB40948),
.ten({ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf1_XU14,ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU14_dbuf0_XU14,ten_measure_currentlimit_XBOTSWZERO,ten_taext_currentlimit_XBOTSWZERO,global_currentlimit_XBOTSWZERO,ten_currentlimit_XBOTSWZERO,global_fetdriver_XBOTSWDRIVER,ten_measure_currentlimit_XBOTSWCURRENT}),
.tma({b0,b0,b0,b1,b0,b1,b0,b1}),
.tmi(tmi[4:0])
);

DFTtm8t dft_hex0x16 (
.G(CELG59462),
.V(CELV96848),
.a({c1,c0}),
.SUB(CELSUB40948),
.ten({noconn_dft_hex0x16_ten_7,ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf1_XU28,ten_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XU28_dbuf0_XU28,ten_currentlimit_delay_XBOTSWZERO_0,ten_currentlimit_delay_XBOTSWZERO_1,ten_currentlimit_delay_XBOTSWZERO_2,ten_currentlimit_delay_XBOTSWZERO_3,ten_currentlimit_delay_XBOTSWZERO_4}),
.tma({c0,c0,c0,c1,c0,c1,c1,c0}),
.tmi(tmi[4:0])
);

drm56 drm_hex0x1c (
.G(CELG59462),
.V(CELV96848),
.d0(e0),
.d1(e1),
.id({e0,e0,e0,e1,e1,e1,e0,e0}),
.SUB(CELSUB40948),
.tmi(tmi[4:0]),
.drm0({noconn_drm56_drm0_7,net_37,net_63,XBOTSWCURRENT_factory_currentlimit_blanking_4,XBOTSWCURRENT_factory_currentlimit_blanking_3,XBOTSWCURRENT_factory_currentlimit_blanking_2,XBOTSWCURRENT_factory_currentlimit_blanking_1,XBOTSWCURRENT_factory_currentlimit_blanking_0}),
.drm1({noconn_drm56_drm1_7,noconn_drm56_drm1_6,noconn_drm56_drm1_5,XBOTSWDRIVER_factory_fetdriver_statusadjust_4,XBOTSWDRIVER_factory_fetdriver_statusadjust_3,XBOTSWDRIVER_factory_fetdriver_statusadjust_2,XBOTSWDRIVER_factory_fetdriver_statusadjust_1,XBOTSWDRIVER_factory_fetdriver_statusadjust_0}),
.drm2({noconn_drm56_drm2_7,noconn_drm56_drm2_6,noconn_drm56_drm2_5,XBOTSWZERO_factory_currentlimit_blanking_4,XBOTSWZERO_factory_currentlimit_blanking_3,XBOTSWZERO_factory_currentlimit_blanking_2,XBOTSWZERO_factory_currentlimit_blanking_1,XBOTSWZERO_factory_currentlimit_blanking_0}),
.drm3({noconn_drm56_drm3_7,noconn_drm56_drm3_6,noconn_drm56_drm3_5,XU11_factory_timingskew_4,XU11_factory_timingskew_3,XU11_factory_timingskew_2,XU11_factory_timingskew_1,XU11_factory_timingskew_0}),
.drm4({noconn_drm56_drm4_7,noconn_drm56_drm4_6,noconn_drm56_drm4_5,XU15_factory_timingskew_4,XU15_factory_timingskew_3,XU15_factory_timingskew_2,XU15_factory_timingskew_1,XU15_factory_timingskew_0}),
.drm5({noconn_drm56_drm5_7,noconn_drm56_drm5_6,noconn_drm56_drm5_5,XU38_factory_timingskew_4,XU38_factory_timingskew_3,XU38_factory_timingskew_2,XU38_factory_timingskew_1,XU38_factory_timingskew_0}),
.drm6({noconn_drm56_drm6_7,noconn_drm56_drm6_6,noconn_drm56_drm6_5,XU41_factory_timingskew_4,XU41_factory_timingskew_3,XU41_factory_timingskew_2,XU41_factory_timingskew_1,XU41_factory_timingskew_0}),
.por0({e0,e1,e1,e0,e0,e0,e0,e0}),
.por1({e0,e0,e0,e0,e0,e0,e0,e0}),
.por2({e0,e0,e0,e0,e0,e0,e0,e0}),
.por3({e0,e0,e0,e0,e0,e1,e1,e0}),
.por4({e0,e0,e0,e0,e1,e0,e0,e0}),
.por5({e0,e0,e0,e0,e0,e1,e1,e0}),
.por6({e0,e0,e0,e0,e0,e1,e1,e0}),
.bypload(e0),
.lastdrm(e0)
);

drm16L drm_hex0x24 (
.G(CELG59462),
.V(CELV96848),
.d0(f0),
.d1(f1),
.id({f0,f0,f1,f0,f0,f1,f0,f0}),
.SUB(CELSUB40948),
.tmi(tmi[4:0]),
.drm0({XBOTSWCURRENT_trim_currentlimit_7,XBOTSWCURRENT_trim_currentlimit_6,XBOTSWCURRENT_trim_currentlimit_5,XBOTSWCURRENT_trim_currentlimit_4,XBOTSWCURRENT_trim_currentlimit_3,XBOTSWCURRENT_trim_currentlimit_2,XBOTSWCURRENT_trim_currentlimit_1,XBOTSWCURRENT_trim_currentlimit_0}),
.drm1({XBOTSWZERO_trim_currentlimit_7,XBOTSWZERO_trim_currentlimit_6,XBOTSWZERO_trim_currentlimit_5,XBOTSWZERO_trim_currentlimit_4,XBOTSWZERO_trim_currentlimit_3,XBOTSWZERO_trim_currentlimit_2,XBOTSWZERO_trim_currentlimit_1,XBOTSWZERO_trim_currentlimit_0}),
.bypload(f0),
.lastdrm(f0)
);

fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWDRIVER XBOTSWDRIVER (
.CELG(CELG59462),
.GATE(net_56),
.HVNEG(PMUDG),
.HVPOS(PMUDV),
.SIMPV(CELV96848),
.fetin(botswon),
.CELSUB(CELSUB40948),
.gate_status(botswstatus),
.global_fetdriver(global_fetdriver_XBOTSWDRIVER),
.enable_fetdriverhv(enable_driver),
.factory_fetdriver_statusadjust({XBOTSWDRIVER_factory_fetdriver_statusadjust_4,XBOTSWDRIVER_factory_fetdriver_statusadjust_3,XBOTSWDRIVER_factory_fetdriver_statusadjust_2,XBOTSWDRIVER_factory_fetdriver_statusadjust_1,XBOTSWDRIVER_factory_fetdriver_statusadjust_0})
);

currentlimitfet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWCURRENT XBOTSWCURRENT (
.IP(IP_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWCURRENT),
.SUB(CELSUB40948),
.CELG(CELG59462),
.SIMPV(MUDV),
.VSENSE(net_112),
.IREPLICA(net_111),
.currentlimit(net_60),
.tdi_currentlimit(tdi_currentlimit_XBOTSWCURRENT),
.ten_currentlimit(ten_currentlimit_XBOTSWCURRENT),
.trim_currentlimit({XBOTSWCURRENT_trim_currentlimit_7,XBOTSWCURRENT_trim_currentlimit_6,XBOTSWCURRENT_trim_currentlimit_5,XBOTSWCURRENT_trim_currentlimit_4,XBOTSWCURRENT_trim_currentlimit_3,XBOTSWCURRENT_trim_currentlimit_2,XBOTSWCURRENT_trim_currentlimit_1,XBOTSWCURRENT_trim_currentlimit_0}),
.TAEXT_CURRENTLIMIT(TAEXT),
.enable_currentlimit(enable_driver),
.global_currentlimit(global_currentlimit_XBOTSWCURRENT),
.measure_currentlimit(botswstatus),
.tdi_currentlimitlive(tdi_currentlimitlive_XBOTSWCURRENT),
.ten_currentlimit_delay({ten_currentlimit_delay_XBOTSWCURRENT_4,ten_currentlimit_delay_XBOTSWCURRENT_3,ten_currentlimit_delay_XBOTSWCURRENT_2,ten_currentlimit_delay_XBOTSWCURRENT_1,ten_currentlimit_delay_XBOTSWCURRENT_0}),
.ten_taext_currentlimit(ten_taext_currentlimit_XBOTSWCURRENT),
.ten_measure_currentlimit(ten_measure_currentlimit_XBOTSWCURRENT),
.factory_currentlimit_blanking({XBOTSWCURRENT_factory_currentlimit_blanking_4,XBOTSWCURRENT_factory_currentlimit_blanking_3,XBOTSWCURRENT_factory_currentlimit_blanking_2,XBOTSWCURRENT_factory_currentlimit_blanking_1,XBOTSWCURRENT_factory_currentlimit_blanking_0})
);

STONEnoconn XNCnoconn_drm56_drm0_7 (
.noconn(noconn_drm56_drm0_7)
);

STONEnoconn XNCnoconn_drm56_drm1_5 (
.noconn(noconn_drm56_drm1_5)
);

STONEnoconn XNCnoconn_drm56_drm1_6 (
.noconn(noconn_drm56_drm1_6)
);

STONEnoconn XNCnoconn_drm56_drm1_7 (
.noconn(noconn_drm56_drm1_7)
);

STONEnoconn XNCnoconn_drm56_drm2_5 (
.noconn(noconn_drm56_drm2_5)
);

STONEnoconn XNCnoconn_drm56_drm2_6 (
.noconn(noconn_drm56_drm2_6)
);

STONEnoconn XNCnoconn_drm56_drm2_7 (
.noconn(noconn_drm56_drm2_7)
);

STONEnoconn XNCnoconn_drm56_drm3_5 (
.noconn(noconn_drm56_drm3_5)
);

STONEnoconn XNCnoconn_drm56_drm3_6 (
.noconn(noconn_drm56_drm3_6)
);

STONEnoconn XNCnoconn_drm56_drm3_7 (
.noconn(noconn_drm56_drm3_7)
);

STONEnoconn XNCnoconn_drm56_drm4_5 (
.noconn(noconn_drm56_drm4_5)
);

STONEnoconn XNCnoconn_drm56_drm4_6 (
.noconn(noconn_drm56_drm4_6)
);

STONEnoconn XNCnoconn_drm56_drm4_7 (
.noconn(noconn_drm56_drm4_7)
);

STONEnoconn XNCnoconn_drm56_drm5_5 (
.noconn(noconn_drm56_drm5_5)
);

STONEnoconn XNCnoconn_drm56_drm5_6 (
.noconn(noconn_drm56_drm5_6)
);

STONEnoconn XNCnoconn_drm56_drm5_7 (
.noconn(noconn_drm56_drm5_7)
);

STONEnoconn XNCnoconn_drm56_drm6_5 (
.noconn(noconn_drm56_drm6_5)
);

STONEnoconn XNCnoconn_drm56_drm6_6 (
.noconn(noconn_drm56_drm6_6)
);

STONEnoconn XNCnoconn_drm56_drm6_7 (
.noconn(noconn_drm56_drm6_7)
);

STONEnoconn XNCnoconn_dft_hex0x16_ten_7 (
.noconn(noconn_dft_hex0x16_ten_7)
);

endmodule

