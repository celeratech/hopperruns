module dftprobe_XLOOP_XCONTROL_XU71 (i,tdi_STEPDOWNalgorithmCONTROL1p3_topstate,ten_STEPDOWNalgorithmCONTROL1p3_topstate,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_topstate;
input  ten_STEPDOWNalgorithmCONTROL1p3_topstate;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

