//Celera:delayfixed_XU1_XSTEPDOWN_XLOOP_XFEEDBACK_XU1_XU4
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:rise
module delayfixed_XU1_XSTEPDOWN_XLOOP_XFEEDBACK_XU1_XU4 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

