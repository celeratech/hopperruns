//Celera:switchtswitch_XLOOP_XREGULATION_XU7_XU10
//Celera Confidential Symbol Generator
//1000 Ohm tswitchSwitch
module switchtswitch_XLOOP_XREGULATION_XU7_XU10 (CELV,O,I,enable_switch,CELG,CELSUB);
input CELV;
input I;
input enable_switch;
inout O;
input CELG;
input CELSUB;
endmodule

