//Celera:delay0_fetdriver_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWDRIVER_Xstatus
//TYPE: fixed 20ns
module delay0_fetdriver_XLOOP_XDRIVER_XBOTDRIVER_XBOTSWDRIVER_Xstatus (i, CELV, o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELSUB;
input CELG;
endmodule

