//Celera:capacitorfixed_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU27
//Celera Confidential Symbol Generator
//CAPACITOR CONTROL:capacitor
//VALUE: 30.00pF TYPE:mim
module capacitorfixed_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU27 (CP,
CN);
inout CP;
inout CN;
endmodule

