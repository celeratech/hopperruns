module dftprobe_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU78 (i,tdi_STEPDOWNalgorithmCONTROL0p2_botstate,ten_STEPDOWNalgorithmCONTROL0p2_botstate,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL0p2_botstate;
input  ten_STEPDOWNalgorithmCONTROL0p2_botstate;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

