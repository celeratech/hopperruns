//Celera:dbuf_XLOOP_XREG_XDEBUG_XU11
//Celera Confidential Symbol Generator
//Digital Buffer
module dbuf_XLOOP_XREG_XDEBUG_XU11 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

