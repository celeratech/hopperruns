module dftprobe_XU1_XSERVICE_XATESERVICE_XU5 (i,tdi_stvbias,ten_stvbias,CELG,CELSUB,CELV);
input  i;
output  tdi_stvbias;
input  ten_stvbias;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

