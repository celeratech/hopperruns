module dftprobe_XLOOP_XREG_XDEBUG_XU2 (i,tdi_REGstartup,ten_REGstartup,CELG,CELSUB,CELV);
input  i;
output  tdi_REGstartup;
input  ten_REGstartup;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

