module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU78 (i,tdi_STEPDOWNalgorithmCORE0p0_FAULT,ten_STEPDOWNalgorithmCORE0p0_FAULT,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_FAULT;
input  ten_STEPDOWNalgorithmCORE0p0_FAULT;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

