//Celera:inv_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU1
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU1 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

