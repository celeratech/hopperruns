//Celera:levelshifter0H2L_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xstatusout
//Celera Confidential Symbol Generator
//Direction: high2low, Maximum high voltage:36V 
//Enable pin:yes
module levelshifter0H2L_fetdriver_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XU9_Xstatusout (SIMPV,CELSUB,HVPOS,HVNEG,in,out,
enable_levelshifter,
CELG);
input SIMPV;
input CELG;
input CELSUB;
input HVPOS;
input HVNEG;
input in;
output out;
input enable_levelshifter;
endmodule

