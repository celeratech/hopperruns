//Celera:resistor_XU1_XSERVICE_XOSCSERVICE_XU4
//Celera Confidential Symbol Generator
//RESISTOR:50.00KOhm TYPE:poly Adjust:25.00Kohm DFT:no
module resistor_XU1_XSERVICE_XOSCSERVICE_XU4 (RP,
CELV,
CELG,
CELSUB,
adjust_resistor,
RN);
inout RP;
inout RN;
input CELV;
input CELG;
input CELSUB;
input [1:0] adjust_resistor;
endmodule

