//Celera:delayfixed_XLOOP_XCONTROL_XU12_XU19
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:both
module delayfixed_XLOOP_XCONTROL_XU12_XU19 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

