//Celera:tie_XLOOP_XCONTROL_XU34_XU31
//Celera Confidential Symbol Generator
//TIE
module tie_XLOOP_XCONTROL_XU34_XU31 (CELV,CELG,a0,SUB);
input CELV;
input CELG;
output a0;
input SUB;
endmodule

