module dftprobe_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU9 (i,tdi_topswipeak,ten_topswipeak,CELG,CELSUB,CELV);
input  i;
output  tdi_topswipeak;
input  ten_topswipeak;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

