module dfthijack_XLOOP_XATE_XU3 (HJendrivero,CELG,CELV,CELSUB,ten_HJendriverenable,ten_HJendriverstatus,HJendriver);
output  HJendrivero;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJendriverenable;
input  ten_HJendriverstatus;
input  HJendriver;
endmodule

