module dftprobe_XLOOP_XDRIVER_XDEBUG_XU18 (i,tdi_DRVbotswzcross,ten_DRVbotswzcross,CELG,CELSUB,CELV);
input  i;
output  tdi_DRVbotswzcross;
input  ten_DRVbotswzcross;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

