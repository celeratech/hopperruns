module dftprobe_XLOOP_XCONTROL_XU65 (i,tdi_STEPDOWNalgorithmCONTROL1p3_FAULT,ten_STEPDOWNalgorithmCONTROL1p3_FAULT,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_FAULT;
input  ten_STEPDOWNalgorithmCONTROL1p3_FAULT;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

