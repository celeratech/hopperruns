module dftprobe_XLOOP_XCONTROL_XU67 (i,tdi_STEPDOWNalgorithmCONTROL1p3_IDLE,ten_STEPDOWNalgorithmCONTROL1p3_IDLE,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_IDLE;
input  ten_STEPDOWNalgorithmCONTROL1p3_IDLE;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

