//Celera:decoder2_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU3_XU2
//Celera Confidential Symbol Generator
//DECODER
module decoder2_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU3_XU2 (CELV,i,o,
CELG,SUB);
input CELV;
input [1:0] i;
output [3:0] o;
input CELG;
input SUB;
endmodule

