// Celera Brick Generator Confidential
//CORE:capacitorfixed
//NAME:capacitorfixed_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU27
//GENERATOR REVISION:0.3.4
//VALUE:30.00Kohms
//Initial Voltage:0V
//TYPE:mim
//VMAX:6V
//DFT:no
//KELVIN:no

//Celera Confidential Do Not Copy mim34_2f30p0x28p9
//Celera Confidential Symbol Generator
//Type mim :30.00pF Capacitor
module mim34_2f30p0x28p9 (CP, CN);
inout CP;
inout CN;
endmodule

//Celera Confidential Do Not Copy capacitorfixed_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU27
//Celera Confidential Symbol Generator
//CAPACITOR CONTROL:capacitor
//VALUE: 30.00pF TYPE:mim
module capacitorfixed_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU2_XU27 (CP,
CN);
inout CP;
inout CN;

//Celera Confidential Do Not Copy Core_
mim34_2f30p0x28p9 XCore_0(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_1(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_2(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_3(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_4(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_5(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_6(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_7(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_8(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_9(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_10(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_11(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_12(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_13(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_14(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_15(
.CP (CP),
.CN (CN)
);
mim34_2f30p0x28p9 XCore_16(
.CP (CP),
.CN (CN)
);

//Celera Confidential Do Not Copy //DieSize,mim34_2f30p0x28p9

//Die Size Calculator mim34_2f30p0x28p9
//,diesize,mim34_2f30p0x28p9,17

//Celera Confidential Do Not Copy Module End
//Celera Schematic Generator
endmodule
