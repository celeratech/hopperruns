module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU89 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_regulation,ten_STEPDOWNalgorithmCORE0p0_enable_regulation,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_enable_regulation;
input  ten_STEPDOWNalgorithmCORE0p0_enable_regulation;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

