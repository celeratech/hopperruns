//Celera:oscillatorcrude_XU1_XSTEPDOWN_XSOFTSTART_XU9_XU9
//Celera Confidential Symbol Generator
//VMAX:globalV,Crude:256.000KHz
module oscillatorcrude_XU1_XSTEPDOWN_XSOFTSTART_XU9_XU9 (SIMPV,ok_oscillator,osc,global_oscillator,
enable_oscillator,
IP,
CELG,SENSE_G,CELSUB);
input SIMPV;
output ok_oscillator;
output osc;
input global_oscillator;
input IP;
input enable_oscillator;
input CELG;
input SENSE_G;
input CELSUB;
endmodule

