//Celera:inv_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU2
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU2 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

