module dftprobe_XU1_XSTEPDOWN_XLOOP_XREGULATION_XU7_XU15 (i,TAI_REGULATIONvc,ten_REGULATIONvc,CELG,CELSUB,CELV);
input  i;
output  TAI_REGULATIONvc;
input  ten_REGULATIONvc;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

