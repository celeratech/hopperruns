module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU84 (i,tdi_STEPDOWNalgorithmCORE0p0_enable_fault,ten_STEPDOWNalgorithmCORE0p0_enable_fault,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_enable_fault;
input  ten_STEPDOWNalgorithmCORE0p0_enable_fault;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

