//Celera:resistordivider_vbuffer_XU1_XSTEPDOWN_XPOWERGOOD_XU3_XU8_Xrfb
//Celera Confidential Symbol Generator
//VMAX:6V R:1000.0KOhm 1Taps
module resistordivider_vbuffer_XU1_XSTEPDOWN_XPOWERGOOD_XU3_XU8_Xrfb (TOP,
TAP0,
CELG, BOTTOM);
inout TOP;
output TAP0;
input CELG;
inout BOTTOM;
endmodule

