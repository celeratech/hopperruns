//Celera:dff_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU9_XU19
//Celera Confidential Symbol Generator
//DFF latch
module dff_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU9_XU19 (CELV,CELG,d,rb,ck,q,qb,SUB );
input CELV;
input CELG;
input d;
input rb;
input ck;
input SUB;
output q;
output qb;
endmodule

