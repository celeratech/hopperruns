//Celera:inv_XLOOP_XDRIVER_XATEDRIVER_XU22_XU15
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XLOOP_XDRIVER_XATEDRIVER_XU22_XU15 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

