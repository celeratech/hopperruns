//Celera:delayfixed_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU15_XU6
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:both
module delayfixed_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU15_XU6 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

