//Celera:comparatorgnd_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU2
//Celera Confidential Symbol Generator
//Threshold: 50 falling
module comparatorgnd_XU1_XSTEPDOWN_XDISCHARGE_XU2_XU3_XU2 (SIMPV,INPUT,out_comparator,IP,
enable_comparator,global_comparator,
sense_CELG,CELSUB,CELG);
input SIMPV;
input INPUT;
output out_comparator;
input IP;
input enable_comparator;
input global_comparator;
input sense_CELG;
input CELG;
input CELSUB;
endmodule

