//Celera:levelshifter0H2L_fetdriver_XLOOP_XDRIVER_XTOPSW_XU12_Xstatusout
//Celera Confidential Symbol Generator
//Direction: high2low, Maximum high voltage:36V 
//Enable pin:yes
module levelshifter0H2L_fetdriver_XLOOP_XDRIVER_XTOPSW_XU12_Xstatusout (SIMPV,CELSUB,HVPOS,HVNEG,in,out,
enable_levelshifter,
CELG);
input SIMPV;
input CELG;
input CELSUB;
input HVPOS;
input HVNEG;
input in;
output out;
input enable_levelshifter;
endmodule

