module dfthijack_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU5 (hjtopstateo,CELG,CELV,CELSUB,ten_hjtopstateenable,ten_hjtopstatestatus,hjtopstate);
output  hjtopstateo;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_hjtopstateenable;
input  ten_hjtopstatestatus;
input  hjtopstate;
endmodule

