//Celera:vbuffer_XU1_XSTEPDOWN_XSOFTSTART_XU8_XU19
//Celera Confidential Symbol Generator
//GAIN:1.1 Input:p with 1000K Impedance
module vbuffer_XU1_XSTEPDOWN_XSOFTSTART_XU8_XU19 (SIMPV,IN,IP,OUT,enable_vbuffer,ok_vbuffer,global_vbuffer,
GNDSENSE,
CELG,CELSUB);
input SIMPV;
input IN;
input IP;
output OUT;
input enable_vbuffer;
output ok_vbuffer;
input global_vbuffer;
input GNDSENSE;
input CELG;
input CELSUB;
endmodule

