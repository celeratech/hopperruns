module dftprobe_XU1_XSTEPDOWN_XLOOP_XDRIVER_XATEDRIVER_XU10 (i,tdi_topswstatus,ten_topswstatus,CELG,CELSUB,CELV);
input  i;
output  tdi_topswstatus;
input  ten_topswstatus;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

