//Celera:feedbackdivider_XLOOP_XFEEDBACK_XFB_XU2
//Celera Confidential Symbol Generator
//Type: control, Feedback Voltage: 1V, Disconnect Pin: pin, P Offset: 0%, N Offset: 0%, Bias Current: 2, DFT: no
//VOUT0:1.2V, VOUT1: 1.5V, VOUT2: 1.8V, VOUT3: 2V, VOUT4: 2.5V, VOUT5: 3.3V, VOUT6: 4.2V, VOUT7: 5V
module feedbackdivider_XLOOP_XFEEDBACK_XFB_XU2 (CELV,SUB,SENSE_FEEDBACKDIVIDER,FEEDBACKDIVIDER_FB,ten,RTN,
pin1,pin2,pin3,
enable_feedbackdivider,
CELG);
input CELV;
input SUB;
input SENSE_FEEDBACKDIVIDER;
output FEEDBACKDIVIDER_FB;
input ten;
input RTN;
input pin1;
input pin2;
input pin3;
input enable_feedbackdivider;
input CELG;
endmodule

