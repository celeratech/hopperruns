module dftprobe_XU1_XSTEPDOWN_XLOOP_XFEEDBACK_XU2_XU2 (i,tdi_FEEDBACKtime,ten_FEEDBACKtime,CELG,CELSUB,CELV);
input  i;
output  tdi_FEEDBACKtime;
input  ten_FEEDBACKtime;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

