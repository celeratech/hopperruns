//Celera:voltage2current_XLOOP_XREGULATION_XU2_XU3
//Celera Confidential Symbol Generator
//Gain: 10, Direction: source, Iout Clamp: no
//DFT:no, Accuracy: no, Input Stage Type: p
module voltage2current_XLOOP_XREGULATION_XU2_XU3 (CELV,SUB,enable_voltage2current,IP,ok_voltage2current,IOUT,VIN,ten,
CELG);
input CELV;
input SUB;
input enable_voltage2current;
input IP;
output ok_voltage2current;
output IOUT;
input VIN;
input ten;
input CELG;
endmodule

