//Celera:srlatch_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU15_XU12
//Celera Confidential Symbol Generator
//SR Latch
module srlatch_XU1_XSTEPDOWN_XLOOP_XCONTROL_XU15_XU12 (CELV,CELG,s,r,rb,q,qb,SUB);
input CELV;
input CELG;
input s;
input r;
input rb;
input SUB;
output q;
output qb;
endmodule

