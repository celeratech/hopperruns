//Celera:levelshifter0H2L_currentlimitfet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XTOPSWCURRENT_Xls
//Celera Confidential Symbol Generator
//Direction: high2low, Maximum high voltage:36V 
//Enable pin:yes
module levelshifter0H2L_currentlimitfet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU6_XTOPSWCURRENT_Xls (SIMPV,CELSUB,HVPOS,HVNEG,in,out,
enable_levelshifter,
CELG);
input SIMPV;
input CELG;
input CELSUB;
input HVPOS;
input HVNEG;
input in;
output out;
input enable_levelshifter;
endmodule

