module dfthijack_XLOOP_XDRIVER_XDEBUG_XU5 (HJdrvtso,CELG,CELV,CELSUB,ten_HJdrvtsenable,ten_HJdrvtsstatus,HJdrvts);
output  HJdrvtso;
input  CELG;
input  CELV;
input  CELSUB;
input  ten_HJdrvtsenable;
input  ten_HJdrvtsstatus;
input  HJdrvts;
endmodule

