module dftprobe_XLOOP_XCONTROL_XU69 (i,tdi_STEPDOWNalgorithmCONTROL1p3_BOTTOM,ten_STEPDOWNalgorithmCONTROL1p3_BOTTOM,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCONTROL1p3_BOTTOM;
input  ten_STEPDOWNalgorithmCONTROL1p3_BOTTOM;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

