//Celera:timingskew_XLOOP_XDRIVER_XBBM_XU14
//Celera Confidential Symbol Generator
//TYPE:rise Bits:5 with 1.0ns LSB
module timingskew_XLOOP_XDRIVER_XBBM_XU14 (CELV,in,out,
factory_timingskew,
CELG,CELSUB);
input CELV;
input in;
output out;
input [4:0] factory_timingskew;
input CELG;
input CELSUB;
endmodule

