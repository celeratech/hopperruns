//Celera:delayfixed_XU1_XSTEPDOWN_XPOWERGOOD_XU13_XU4
//Celera Confidential Symbol Generator
//TYPE:fixed Egde:fall
module delayfixed_XU1_XSTEPDOWN_XPOWERGOOD_XU13_XU4 (CELV,i,o,
CELG,CELSUB);
input CELV;
input i;
output o;
input CELG;
input CELSUB;
endmodule

