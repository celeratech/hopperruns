//Celera:srlatch_XLOOP_XCONTROL_XU32_XU13
//Celera Confidential Symbol Generator
//SR Latch
module srlatch_XLOOP_XCONTROL_XU32_XU13 (CELV,CELG,s,r,rb,q,qb,SUB);
input CELV;
input CELG;
input s;
input r;
input rb;
input SUB;
output q;
output qb;
endmodule

