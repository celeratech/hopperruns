//Celera:inv_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU23_XU5
//Celera Confidential Symbol Generator
//5V Inverter
module inv_XU1_XSTEPDOWN_XSOFTSTART_XU1_XU23_XU5 (CELV,CELG,i,o,SUB);
input CELV;
input CELG;
input i;
input SUB;
output o;
endmodule

