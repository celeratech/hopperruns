//Celera:fetdriver_XLOOP_XDRIVER_XTOPDRIVER_XTOPSWDRIVER
//Celera Confidential Symbol Generator
//FET DRIVER 'n' Type 4 Ron 2 Roff 
//Input 36V Levelshifter
//Gate Sense None
//DFT no
module fetdriver_XLOOP_XDRIVER_XTOPDRIVER_XTOPSWDRIVER (HVPOS,enable_fetdriverhv,global_fetdriver,fetin,GATE,gate_status,
CELG,
SIMPV,
enable_fetdriver,
HVNEG,CELSUB); 
input HVPOS;
input enable_fetdriverhv;
input global_fetdriver;
input fetin;
output GATE;
output gate_status;
input SIMPV;
input CELG;
input enable_fetdriver;
input HVNEG;
input CELSUB;
endmodule

