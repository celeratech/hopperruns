module dftprobe_XU1_XSTEPDOWN_XCORESTATE_XU80 (i,tdi_STEPDOWNalgorithmCORE0p0_POWERDOWN,ten_STEPDOWNalgorithmCORE0p0_POWERDOWN,CELG,CELSUB,CELV);
input  i;
output  tdi_STEPDOWNalgorithmCORE0p0_POWERDOWN;
input  ten_STEPDOWNalgorithmCORE0p0_POWERDOWN;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

