module dftprobe_XLOOP_XDRIVER_XDEBUG_XU20 (i,tdi_DRVSLOPETRIM,ten_DRVSLOPETRIM,CELG,CELSUB,CELV);
input  i;
output  tdi_DRVSLOPETRIM;
input  ten_DRVSLOPETRIM;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

