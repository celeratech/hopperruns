//Celera:fet_fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZREP_Xfet
//Celera Confidential Symbol Generator
//power NMOS:Ron:0.200 Ohm
//Vgs 6V Vds 30V
//Kelvin:no

module fet_fet_XU1_XSTEPDOWN_XLOOP_XDRIVER_XU2_XBOTSWZREP_Xfet (GATE,SOURCE,DRAIN,SUB);
input GATE;
inout SOURCE;
inout DRAIN;
input SUB;
endmodule

