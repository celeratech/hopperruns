module dftprobe_XU1_XSTEPDOWN_XFAULT_XU1_XU13 (i,tdi_FAULTtime,ten_FAULTtime,CELG,CELSUB,CELV);
input  i;
output  tdi_FAULTtime;
input  ten_FAULTtime;
input  CELG;
input  CELSUB;
input  CELV;
endmodule

